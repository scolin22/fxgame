// nios_system.v

// Generated using ACDS version 12.0sp2 263 at 2014.01.19.20:59:23

`timescale 1 ps / 1 ps
module nios_system (
		input  wire [7:0]  switches_export,      //       switches.export
		output wire [7:0]  leds_export,          //           leds.export
		inout  wire [15:0] sram_DQ,              //           sram.DQ
		output wire [17:0] sram_ADDR,            //               .ADDR
		output wire        sram_LB_N,            //               .LB_N
		output wire        sram_UB_N,            //               .UB_N
		output wire        sram_CE_N,            //               .CE_N
		output wire        sram_OE_N,            //               .OE_N
		output wire        sram_WE_N,            //               .WE_N
		output wire [11:0] sdram_wire_addr,      //     sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,        //               .ba
		output wire        sdram_wire_cas_n,     //               .cas_n
		output wire        sdram_wire_cke,       //               .cke
		output wire        sdram_wire_cs_n,      //               .cs_n
		inout  wire [15:0] sdram_wire_dq,        //               .dq
		output wire [1:0]  sdram_wire_dqm,       //               .dqm
		output wire        sdram_wire_ras_n,     //               .ras_n
		output wire        sdram_wire_we_n,      //               .we_n
		input  wire        reset_reset_n,        //          reset.reset_n
		output wire        vga_controller_CLK,   // vga_controller.CLK
		output wire        vga_controller_HS,    //               .HS
		output wire        vga_controller_VS,    //               .VS
		output wire        vga_controller_BLANK, //               .BLANK
		output wire        vga_controller_SYNC,  //               .SYNC
		output wire [9:0]  vga_controller_R,     //               .R
		output wire [9:0]  vga_controller_G,     //               .G
		output wire [9:0]  vga_controller_B,     //               .B
		input  wire        clk_clk,              //            clk.clk
		output wire        sdram_clk_clk,        //      sdram_clk.clk
		inout  wire [7:0]  lcd_data_DATA,        //       lcd_data.DATA
		output wire        lcd_data_ON,          //               .ON
		output wire        lcd_data_BLON,        //               .BLON
		output wire        lcd_data_EN,          //               .EN
		output wire        lcd_data_RS,          //               .RS
		output wire        lcd_data_RW           //               .RW
	);

	wire          clocks_sys_clk_clk;                                                                                         // clocks:sys_clk -> [LEDs:clk, LEDs_s1_translator:clk, LEDs_s1_translator_avalon_universal_slave_0_agent:clk, LEDs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, addr_router:clk, addr_router_001:clk, addr_router_002:clk, alpha_blender:clk, burst_adapter:clk, burst_adapter_001:clk, burst_adapter_002:clk, burst_adapter_003:clk, char_drawer:clk, char_drawer_avalon_char_buffer_slave_translator:clk, char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:clk, char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, char_drawer_avalon_char_control_slave_translator:clk, char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:clk, char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, character_lcd_0:clk, character_lcd_0_avalon_lcd_slave_translator:clk, character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:clk, character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, cmd_xbar_demux:clk, cmd_xbar_demux_001:clk, cmd_xbar_demux_002:clk, cmd_xbar_mux:clk, cmd_xbar_mux_001:clk, cmd_xbar_mux_002:clk, cmd_xbar_mux_007:clk, id_router:clk, id_router_001:clk, id_router_002:clk, id_router_003:clk, id_router_004:clk, id_router_005:clk, id_router_006:clk, id_router_007:clk, id_router_008:clk, id_router_009:clk, id_router_010:clk, irq_mapper:clk, jtag_uart_0:clk, jtag_uart_0_avalon_jtag_slave_translator:clk, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:clk, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, limiter:clk, nios2_processor:clk, nios2_processor_data_master_translator:clk, nios2_processor_data_master_translator_avalon_universal_master_0_agent:clk, nios2_processor_instruction_master_translator:clk, nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:clk, nios2_processor_jtag_debug_module_translator:clk, nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:clk, nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, onchip_memory2_0:clk, onchip_memory2_0_s1_translator:clk, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:clk, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pixel_buffer:clk, pixel_buffer_avalon_sram_slave_translator:clk, pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:clk, pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pixel_buffer_dma:clk, pixel_buffer_dma_avalon_control_slave_translator:clk, pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:clk, pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pixel_buffer_dma_avalon_pixel_dma_master_translator:clk, pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:clk, rgb_resampler:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_002:clk, rsp_xbar_demux_003:clk, rsp_xbar_demux_004:clk, rsp_xbar_demux_005:clk, rsp_xbar_demux_006:clk, rsp_xbar_demux_007:clk, rsp_xbar_demux_008:clk, rsp_xbar_demux_009:clk, rsp_xbar_demux_010:clk, rsp_xbar_mux:clk, rsp_xbar_mux_001:clk, rst_controller:clk, scaler:clk, sdram:clk, sdram_s1_translator:clk, sdram_s1_translator_avalon_universal_slave_0_agent:clk, sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, switches:clk, switches_s1_translator:clk, switches_s1_translator_avalon_universal_slave_0_agent:clk, switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, video_fifo:clk_stream_in, width_adapter:clk, width_adapter_001:clk, width_adapter_002:clk, width_adapter_003:clk, width_adapter_004:clk, width_adapter_005:clk, width_adapter_006:clk, width_adapter_007:clk, width_adapter_008:clk, width_adapter_009:clk]
	wire          pixel_buffer_dma_avalon_pixel_source_endofpacket;                                                           // pixel_buffer_dma:stream_endofpacket -> rgb_resampler:stream_in_endofpacket
	wire          pixel_buffer_dma_avalon_pixel_source_valid;                                                                 // pixel_buffer_dma:stream_valid -> rgb_resampler:stream_in_valid
	wire          pixel_buffer_dma_avalon_pixel_source_startofpacket;                                                         // pixel_buffer_dma:stream_startofpacket -> rgb_resampler:stream_in_startofpacket
	wire   [15:0] pixel_buffer_dma_avalon_pixel_source_data;                                                                  // pixel_buffer_dma:stream_data -> rgb_resampler:stream_in_data
	wire          pixel_buffer_dma_avalon_pixel_source_ready;                                                                 // rgb_resampler:stream_in_ready -> pixel_buffer_dma:stream_ready
	wire          rgb_resampler_avalon_rgb_source_endofpacket;                                                                // rgb_resampler:stream_out_endofpacket -> scaler:stream_in_endofpacket
	wire          rgb_resampler_avalon_rgb_source_valid;                                                                      // rgb_resampler:stream_out_valid -> scaler:stream_in_valid
	wire          rgb_resampler_avalon_rgb_source_startofpacket;                                                              // rgb_resampler:stream_out_startofpacket -> scaler:stream_in_startofpacket
	wire   [29:0] rgb_resampler_avalon_rgb_source_data;                                                                       // rgb_resampler:stream_out_data -> scaler:stream_in_data
	wire          rgb_resampler_avalon_rgb_source_ready;                                                                      // scaler:stream_in_ready -> rgb_resampler:stream_out_ready
	wire          clocks_vga_clk_clk;                                                                                         // clocks:VGA_CLK -> [rst_controller_002:clk, vga_controller:clk, video_fifo:clk_stream_out]
	wire          video_fifo_avalon_dc_buffer_source_endofpacket;                                                             // video_fifo:stream_out_endofpacket -> vga_controller:endofpacket
	wire          video_fifo_avalon_dc_buffer_source_valid;                                                                   // video_fifo:stream_out_valid -> vga_controller:valid
	wire          video_fifo_avalon_dc_buffer_source_startofpacket;                                                           // video_fifo:stream_out_startofpacket -> vga_controller:startofpacket
	wire   [29:0] video_fifo_avalon_dc_buffer_source_data;                                                                    // video_fifo:stream_out_data -> vga_controller:data
	wire          video_fifo_avalon_dc_buffer_source_ready;                                                                   // vga_controller:ready -> video_fifo:stream_out_ready
	wire          char_drawer_avalon_char_source_endofpacket;                                                                 // char_drawer:stream_endofpacket -> alpha_blender:foreground_endofpacket
	wire          char_drawer_avalon_char_source_valid;                                                                       // char_drawer:stream_valid -> alpha_blender:foreground_valid
	wire          char_drawer_avalon_char_source_startofpacket;                                                               // char_drawer:stream_startofpacket -> alpha_blender:foreground_startofpacket
	wire   [39:0] char_drawer_avalon_char_source_data;                                                                        // char_drawer:stream_data -> alpha_blender:foreground_data
	wire          char_drawer_avalon_char_source_ready;                                                                       // alpha_blender:foreground_ready -> char_drawer:stream_ready
	wire          scaler_avalon_scaler_source_endofpacket;                                                                    // scaler:stream_out_endofpacket -> alpha_blender:background_endofpacket
	wire          scaler_avalon_scaler_source_valid;                                                                          // scaler:stream_out_valid -> alpha_blender:background_valid
	wire          scaler_avalon_scaler_source_startofpacket;                                                                  // scaler:stream_out_startofpacket -> alpha_blender:background_startofpacket
	wire   [29:0] scaler_avalon_scaler_source_data;                                                                           // scaler:stream_out_data -> alpha_blender:background_data
	wire          scaler_avalon_scaler_source_ready;                                                                          // alpha_blender:background_ready -> scaler:stream_out_ready
	wire          alpha_blender_avalon_blended_source_endofpacket;                                                            // alpha_blender:output_endofpacket -> video_fifo:stream_in_endofpacket
	wire          alpha_blender_avalon_blended_source_valid;                                                                  // alpha_blender:output_valid -> video_fifo:stream_in_valid
	wire          alpha_blender_avalon_blended_source_startofpacket;                                                          // alpha_blender:output_startofpacket -> video_fifo:stream_in_startofpacket
	wire   [29:0] alpha_blender_avalon_blended_source_data;                                                                   // alpha_blender:output_data -> video_fifo:stream_in_data
	wire          alpha_blender_avalon_blended_source_ready;                                                                  // video_fifo:stream_in_ready -> alpha_blender:output_ready
	wire          nios2_processor_instruction_master_waitrequest;                                                             // nios2_processor_instruction_master_translator:av_waitrequest -> nios2_processor:i_waitrequest
	wire   [24:0] nios2_processor_instruction_master_address;                                                                 // nios2_processor:i_address -> nios2_processor_instruction_master_translator:av_address
	wire          nios2_processor_instruction_master_read;                                                                    // nios2_processor:i_read -> nios2_processor_instruction_master_translator:av_read
	wire   [31:0] nios2_processor_instruction_master_readdata;                                                                // nios2_processor_instruction_master_translator:av_readdata -> nios2_processor:i_readdata
	wire          nios2_processor_instruction_master_readdatavalid;                                                           // nios2_processor_instruction_master_translator:av_readdatavalid -> nios2_processor:i_readdatavalid
	wire          nios2_processor_data_master_waitrequest;                                                                    // nios2_processor_data_master_translator:av_waitrequest -> nios2_processor:d_waitrequest
	wire   [31:0] nios2_processor_data_master_writedata;                                                                      // nios2_processor:d_writedata -> nios2_processor_data_master_translator:av_writedata
	wire   [24:0] nios2_processor_data_master_address;                                                                        // nios2_processor:d_address -> nios2_processor_data_master_translator:av_address
	wire          nios2_processor_data_master_write;                                                                          // nios2_processor:d_write -> nios2_processor_data_master_translator:av_write
	wire          nios2_processor_data_master_read;                                                                           // nios2_processor:d_read -> nios2_processor_data_master_translator:av_read
	wire   [31:0] nios2_processor_data_master_readdata;                                                                       // nios2_processor_data_master_translator:av_readdata -> nios2_processor:d_readdata
	wire          nios2_processor_data_master_debugaccess;                                                                    // nios2_processor:jtag_debug_module_debugaccess_to_roms -> nios2_processor_data_master_translator:av_debugaccess
	wire    [3:0] nios2_processor_data_master_byteenable;                                                                     // nios2_processor:d_byteenable -> nios2_processor_data_master_translator:av_byteenable
	wire          pixel_buffer_dma_avalon_pixel_dma_master_waitrequest;                                                       // pixel_buffer_dma_avalon_pixel_dma_master_translator:av_waitrequest -> pixel_buffer_dma:master_waitrequest
	wire   [31:0] pixel_buffer_dma_avalon_pixel_dma_master_address;                                                           // pixel_buffer_dma:master_address -> pixel_buffer_dma_avalon_pixel_dma_master_translator:av_address
	wire          pixel_buffer_dma_avalon_pixel_dma_master_lock;                                                              // pixel_buffer_dma:master_arbiterlock -> pixel_buffer_dma_avalon_pixel_dma_master_translator:av_lock
	wire          pixel_buffer_dma_avalon_pixel_dma_master_read;                                                              // pixel_buffer_dma:master_read -> pixel_buffer_dma_avalon_pixel_dma_master_translator:av_read
	wire   [15:0] pixel_buffer_dma_avalon_pixel_dma_master_readdata;                                                          // pixel_buffer_dma_avalon_pixel_dma_master_translator:av_readdata -> pixel_buffer_dma:master_readdata
	wire          pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid;                                                     // pixel_buffer_dma_avalon_pixel_dma_master_translator:av_readdatavalid -> pixel_buffer_dma:master_readdatavalid
	wire   [31:0] nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                 // nios2_processor_jtag_debug_module_translator:av_writedata -> nios2_processor:jtag_debug_module_writedata
	wire    [8:0] nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_address;                                   // nios2_processor_jtag_debug_module_translator:av_address -> nios2_processor:jtag_debug_module_address
	wire          nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                                // nios2_processor_jtag_debug_module_translator:av_chipselect -> nios2_processor:jtag_debug_module_select
	wire          nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_write;                                     // nios2_processor_jtag_debug_module_translator:av_write -> nios2_processor:jtag_debug_module_write
	wire   [31:0] nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                  // nios2_processor:jtag_debug_module_readdata -> nios2_processor_jtag_debug_module_translator:av_readdata
	wire          nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                             // nios2_processor_jtag_debug_module_translator:av_begintransfer -> nios2_processor:jtag_debug_module_begintransfer
	wire          nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                               // nios2_processor_jtag_debug_module_translator:av_debugaccess -> nios2_processor:jtag_debug_module_debugaccess
	wire    [3:0] nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                // nios2_processor_jtag_debug_module_translator:av_byteenable -> nios2_processor:jtag_debug_module_byteenable
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata;                                               // onchip_memory2_0_s1_translator:av_writedata -> onchip_memory2_0:writedata
	wire    [9:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_address;                                                 // onchip_memory2_0_s1_translator:av_address -> onchip_memory2_0:address
	wire          onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect;                                              // onchip_memory2_0_s1_translator:av_chipselect -> onchip_memory2_0:chipselect
	wire          onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken;                                                   // onchip_memory2_0_s1_translator:av_clken -> onchip_memory2_0:clken
	wire          onchip_memory2_0_s1_translator_avalon_anti_slave_0_write;                                                   // onchip_memory2_0_s1_translator:av_write -> onchip_memory2_0:write
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata;                                                // onchip_memory2_0:readdata -> onchip_memory2_0_s1_translator:av_readdata
	wire    [3:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable;                                              // onchip_memory2_0_s1_translator:av_byteenable -> onchip_memory2_0:byteenable
	wire          sdram_s1_translator_avalon_anti_slave_0_waitrequest;                                                        // sdram:za_waitrequest -> sdram_s1_translator:av_waitrequest
	wire   [15:0] sdram_s1_translator_avalon_anti_slave_0_writedata;                                                          // sdram_s1_translator:av_writedata -> sdram:az_data
	wire   [21:0] sdram_s1_translator_avalon_anti_slave_0_address;                                                            // sdram_s1_translator:av_address -> sdram:az_addr
	wire          sdram_s1_translator_avalon_anti_slave_0_chipselect;                                                         // sdram_s1_translator:av_chipselect -> sdram:az_cs
	wire          sdram_s1_translator_avalon_anti_slave_0_write;                                                              // sdram_s1_translator:av_write -> sdram:az_wr_n
	wire          sdram_s1_translator_avalon_anti_slave_0_read;                                                               // sdram_s1_translator:av_read -> sdram:az_rd_n
	wire   [15:0] sdram_s1_translator_avalon_anti_slave_0_readdata;                                                           // sdram:za_data -> sdram_s1_translator:av_readdata
	wire          sdram_s1_translator_avalon_anti_slave_0_readdatavalid;                                                      // sdram:za_valid -> sdram_s1_translator:av_readdatavalid
	wire    [1:0] sdram_s1_translator_avalon_anti_slave_0_byteenable;                                                         // sdram_s1_translator:av_byteenable -> sdram:az_be_n
	wire   [31:0] leds_s1_translator_avalon_anti_slave_0_writedata;                                                           // LEDs_s1_translator:av_writedata -> LEDs:writedata
	wire    [1:0] leds_s1_translator_avalon_anti_slave_0_address;                                                             // LEDs_s1_translator:av_address -> LEDs:address
	wire          leds_s1_translator_avalon_anti_slave_0_chipselect;                                                          // LEDs_s1_translator:av_chipselect -> LEDs:chipselect
	wire          leds_s1_translator_avalon_anti_slave_0_write;                                                               // LEDs_s1_translator:av_write -> LEDs:write_n
	wire   [31:0] leds_s1_translator_avalon_anti_slave_0_readdata;                                                            // LEDs:readdata -> LEDs_s1_translator:av_readdata
	wire    [1:0] switches_s1_translator_avalon_anti_slave_0_address;                                                         // switches_s1_translator:av_address -> switches:address
	wire   [31:0] switches_s1_translator_avalon_anti_slave_0_readdata;                                                        // switches:readdata -> switches_s1_translator:av_readdata
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                                   // jtag_uart_0:av_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                                     // jtag_uart_0_avalon_jtag_slave_translator:av_writedata -> jtag_uart_0:av_writedata
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                       // jtag_uart_0_avalon_jtag_slave_translator:av_address -> jtag_uart_0:av_address
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                                    // jtag_uart_0_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_0:av_chipselect
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                         // jtag_uart_0_avalon_jtag_slave_translator:av_write -> jtag_uart_0:av_write_n
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                          // jtag_uart_0_avalon_jtag_slave_translator:av_read -> jtag_uart_0:av_read_n
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                                      // jtag_uart_0:av_readdata -> jtag_uart_0_avalon_jtag_slave_translator:av_readdata
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_waitrequest;                                // character_lcd_0:waitrequest -> character_lcd_0_avalon_lcd_slave_translator:av_waitrequest
	wire    [7:0] character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_writedata;                                  // character_lcd_0_avalon_lcd_slave_translator:av_writedata -> character_lcd_0:writedata
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_address;                                    // character_lcd_0_avalon_lcd_slave_translator:av_address -> character_lcd_0:address
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_chipselect;                                 // character_lcd_0_avalon_lcd_slave_translator:av_chipselect -> character_lcd_0:chipselect
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_write;                                      // character_lcd_0_avalon_lcd_slave_translator:av_write -> character_lcd_0:write
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_read;                                       // character_lcd_0_avalon_lcd_slave_translator:av_read -> character_lcd_0:read
	wire    [7:0] character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_readdata;                                   // character_lcd_0:readdata -> character_lcd_0_avalon_lcd_slave_translator:av_readdata
	wire   [15:0] pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_writedata;                                    // pixel_buffer_avalon_sram_slave_translator:av_writedata -> pixel_buffer:writedata
	wire   [17:0] pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_address;                                      // pixel_buffer_avalon_sram_slave_translator:av_address -> pixel_buffer:address
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_write;                                        // pixel_buffer_avalon_sram_slave_translator:av_write -> pixel_buffer:write
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_read;                                         // pixel_buffer_avalon_sram_slave_translator:av_read -> pixel_buffer:read
	wire   [15:0] pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdata;                                     // pixel_buffer:readdata -> pixel_buffer_avalon_sram_slave_translator:av_readdata
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid;                                // pixel_buffer:readdatavalid -> pixel_buffer_avalon_sram_slave_translator:av_readdatavalid
	wire    [1:0] pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable;                                   // pixel_buffer_avalon_sram_slave_translator:av_byteenable -> pixel_buffer:byteenable
	wire   [31:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_writedata;                             // pixel_buffer_dma_avalon_control_slave_translator:av_writedata -> pixel_buffer_dma:slave_writedata
	wire    [1:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_address;                               // pixel_buffer_dma_avalon_control_slave_translator:av_address -> pixel_buffer_dma:slave_address
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_write;                                 // pixel_buffer_dma_avalon_control_slave_translator:av_write -> pixel_buffer_dma:slave_write
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_read;                                  // pixel_buffer_dma_avalon_control_slave_translator:av_read -> pixel_buffer_dma:slave_read
	wire   [31:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_readdata;                              // pixel_buffer_dma:slave_readdata -> pixel_buffer_dma_avalon_control_slave_translator:av_readdata
	wire    [3:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_byteenable;                            // pixel_buffer_dma_avalon_control_slave_translator:av_byteenable -> pixel_buffer_dma:slave_byteenable
	wire   [31:0] char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_writedata;                             // char_drawer_avalon_char_control_slave_translator:av_writedata -> char_drawer:ctrl_writedata
	wire          char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_address;                               // char_drawer_avalon_char_control_slave_translator:av_address -> char_drawer:ctrl_address
	wire          char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_chipselect;                            // char_drawer_avalon_char_control_slave_translator:av_chipselect -> char_drawer:ctrl_chipselect
	wire          char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_write;                                 // char_drawer_avalon_char_control_slave_translator:av_write -> char_drawer:ctrl_write
	wire          char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_read;                                  // char_drawer_avalon_char_control_slave_translator:av_read -> char_drawer:ctrl_read
	wire   [31:0] char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_readdata;                              // char_drawer:ctrl_readdata -> char_drawer_avalon_char_control_slave_translator:av_readdata
	wire    [3:0] char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_byteenable;                            // char_drawer_avalon_char_control_slave_translator:av_byteenable -> char_drawer:ctrl_byteenable
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_waitrequest;                            // char_drawer:buf_waitrequest -> char_drawer_avalon_char_buffer_slave_translator:av_waitrequest
	wire    [7:0] char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_writedata;                              // char_drawer_avalon_char_buffer_slave_translator:av_writedata -> char_drawer:buf_writedata
	wire   [12:0] char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_address;                                // char_drawer_avalon_char_buffer_slave_translator:av_address -> char_drawer:buf_address
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_chipselect;                             // char_drawer_avalon_char_buffer_slave_translator:av_chipselect -> char_drawer:buf_chipselect
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_write;                                  // char_drawer_avalon_char_buffer_slave_translator:av_write -> char_drawer:buf_write
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_read;                                   // char_drawer_avalon_char_buffer_slave_translator:av_read -> char_drawer:buf_read
	wire    [7:0] char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_readdata;                               // char_drawer:buf_readdata -> char_drawer_avalon_char_buffer_slave_translator:av_readdata
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_byteenable;                             // char_drawer_avalon_char_buffer_slave_translator:av_byteenable -> char_drawer:buf_byteenable
	wire          nios2_processor_instruction_master_translator_avalon_universal_master_0_waitrequest;                        // nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_processor_instruction_master_translator:uav_waitrequest
	wire    [2:0] nios2_processor_instruction_master_translator_avalon_universal_master_0_burstcount;                         // nios2_processor_instruction_master_translator:uav_burstcount -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] nios2_processor_instruction_master_translator_avalon_universal_master_0_writedata;                          // nios2_processor_instruction_master_translator:uav_writedata -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] nios2_processor_instruction_master_translator_avalon_universal_master_0_address;                            // nios2_processor_instruction_master_translator:uav_address -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          nios2_processor_instruction_master_translator_avalon_universal_master_0_lock;                               // nios2_processor_instruction_master_translator:uav_lock -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          nios2_processor_instruction_master_translator_avalon_universal_master_0_write;                              // nios2_processor_instruction_master_translator:uav_write -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          nios2_processor_instruction_master_translator_avalon_universal_master_0_read;                               // nios2_processor_instruction_master_translator:uav_read -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] nios2_processor_instruction_master_translator_avalon_universal_master_0_readdata;                           // nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_processor_instruction_master_translator:uav_readdata
	wire          nios2_processor_instruction_master_translator_avalon_universal_master_0_debugaccess;                        // nios2_processor_instruction_master_translator:uav_debugaccess -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] nios2_processor_instruction_master_translator_avalon_universal_master_0_byteenable;                         // nios2_processor_instruction_master_translator:uav_byteenable -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          nios2_processor_instruction_master_translator_avalon_universal_master_0_readdatavalid;                      // nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_processor_instruction_master_translator:uav_readdatavalid
	wire          nios2_processor_data_master_translator_avalon_universal_master_0_waitrequest;                               // nios2_processor_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_processor_data_master_translator:uav_waitrequest
	wire    [2:0] nios2_processor_data_master_translator_avalon_universal_master_0_burstcount;                                // nios2_processor_data_master_translator:uav_burstcount -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] nios2_processor_data_master_translator_avalon_universal_master_0_writedata;                                 // nios2_processor_data_master_translator:uav_writedata -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] nios2_processor_data_master_translator_avalon_universal_master_0_address;                                   // nios2_processor_data_master_translator:uav_address -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          nios2_processor_data_master_translator_avalon_universal_master_0_lock;                                      // nios2_processor_data_master_translator:uav_lock -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          nios2_processor_data_master_translator_avalon_universal_master_0_write;                                     // nios2_processor_data_master_translator:uav_write -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          nios2_processor_data_master_translator_avalon_universal_master_0_read;                                      // nios2_processor_data_master_translator:uav_read -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] nios2_processor_data_master_translator_avalon_universal_master_0_readdata;                                  // nios2_processor_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_processor_data_master_translator:uav_readdata
	wire          nios2_processor_data_master_translator_avalon_universal_master_0_debugaccess;                               // nios2_processor_data_master_translator:uav_debugaccess -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] nios2_processor_data_master_translator_avalon_universal_master_0_byteenable;                                // nios2_processor_data_master_translator:uav_byteenable -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          nios2_processor_data_master_translator_avalon_universal_master_0_readdatavalid;                             // nios2_processor_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_processor_data_master_translator:uav_readdatavalid
	wire          pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_waitrequest;                  // pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_waitrequest -> pixel_buffer_dma_avalon_pixel_dma_master_translator:uav_waitrequest
	wire    [1:0] pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_burstcount;                   // pixel_buffer_dma_avalon_pixel_dma_master_translator:uav_burstcount -> pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [15:0] pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_writedata;                    // pixel_buffer_dma_avalon_pixel_dma_master_translator:uav_writedata -> pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_address;                      // pixel_buffer_dma_avalon_pixel_dma_master_translator:uav_address -> pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_address
	wire          pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_lock;                         // pixel_buffer_dma_avalon_pixel_dma_master_translator:uav_lock -> pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_lock
	wire          pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_write;                        // pixel_buffer_dma_avalon_pixel_dma_master_translator:uav_write -> pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_write
	wire          pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_read;                         // pixel_buffer_dma_avalon_pixel_dma_master_translator:uav_read -> pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_read
	wire   [15:0] pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdata;                     // pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_readdata -> pixel_buffer_dma_avalon_pixel_dma_master_translator:uav_readdata
	wire          pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_debugaccess;                  // pixel_buffer_dma_avalon_pixel_dma_master_translator:uav_debugaccess -> pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [1:0] pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_byteenable;                   // pixel_buffer_dma_avalon_pixel_dma_master_translator:uav_byteenable -> pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdatavalid;                // pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> pixel_buffer_dma_avalon_pixel_dma_master_translator:uav_readdatavalid
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                 // nios2_processor_jtag_debug_module_translator:uav_waitrequest -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                  // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios2_processor_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                   // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios2_processor_jtag_debug_module_translator:uav_writedata
	wire   [31:0] nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                     // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios2_processor_jtag_debug_module_translator:uav_address
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                       // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios2_processor_jtag_debug_module_translator:uav_write
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                        // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios2_processor_jtag_debug_module_translator:uav_lock
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                        // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios2_processor_jtag_debug_module_translator:uav_read
	wire   [31:0] nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                    // nios2_processor_jtag_debug_module_translator:uav_readdata -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;               // nios2_processor_jtag_debug_module_translator:uav_readdatavalid -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                 // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios2_processor_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                  // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios2_processor_jtag_debug_module_translator:uav_byteenable
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;          // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;        // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [105:0] nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                 // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;       // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;             // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;     // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [105:0] nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;              // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;             // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;           // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;            // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;           // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // onchip_memory2_0_s1_translator:uav_waitrequest -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> onchip_memory2_0_s1_translator:uav_burstcount
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> onchip_memory2_0_s1_translator:uav_writedata
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                   // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> onchip_memory2_0_s1_translator:uav_address
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                     // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> onchip_memory2_0_s1_translator:uav_write
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                      // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> onchip_memory2_0_s1_translator:uav_lock
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                      // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> onchip_memory2_0_s1_translator:uav_read
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // onchip_memory2_0_s1_translator:uav_readdata -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // onchip_memory2_0_s1_translator:uav_readdatavalid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> onchip_memory2_0_s1_translator:uav_debugaccess
	wire    [3:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> onchip_memory2_0_s1_translator:uav_byteenable
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [105:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                               // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [105:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                          // sdram_s1_translator:uav_waitrequest -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                           // sdram_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdram_s1_translator:uav_burstcount
	wire   [15:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                            // sdram_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sdram_s1_translator:uav_writedata
	wire   [31:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_address;                                              // sdram_s1_translator_avalon_universal_slave_0_agent:m0_address -> sdram_s1_translator:uav_address
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                // sdram_s1_translator_avalon_universal_slave_0_agent:m0_write -> sdram_s1_translator:uav_write
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                 // sdram_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sdram_s1_translator:uav_lock
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                 // sdram_s1_translator_avalon_universal_slave_0_agent:m0_read -> sdram_s1_translator:uav_read
	wire   [15:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                             // sdram_s1_translator:uav_readdata -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                        // sdram_s1_translator:uav_readdatavalid -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                          // sdram_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdram_s1_translator:uav_debugaccess
	wire    [1:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                           // sdram_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdram_s1_translator:uav_byteenable
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                   // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                         // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                 // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [87:0] sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                          // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                         // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                      // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                              // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [87:0] sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                       // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                      // sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                    // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [15:0] sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                     // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                    // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                           // LEDs_s1_translator:uav_waitrequest -> LEDs_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                            // LEDs_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> LEDs_s1_translator:uav_burstcount
	wire   [31:0] leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                             // LEDs_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> LEDs_s1_translator:uav_writedata
	wire   [31:0] leds_s1_translator_avalon_universal_slave_0_agent_m0_address;                                               // LEDs_s1_translator_avalon_universal_slave_0_agent:m0_address -> LEDs_s1_translator:uav_address
	wire          leds_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                 // LEDs_s1_translator_avalon_universal_slave_0_agent:m0_write -> LEDs_s1_translator:uav_write
	wire          leds_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                  // LEDs_s1_translator_avalon_universal_slave_0_agent:m0_lock -> LEDs_s1_translator:uav_lock
	wire          leds_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                  // LEDs_s1_translator_avalon_universal_slave_0_agent:m0_read -> LEDs_s1_translator:uav_read
	wire   [31:0] leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                              // LEDs_s1_translator:uav_readdata -> LEDs_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                         // LEDs_s1_translator:uav_readdatavalid -> LEDs_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                           // LEDs_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> LEDs_s1_translator:uav_debugaccess
	wire    [3:0] leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                            // LEDs_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> LEDs_s1_translator:uav_byteenable
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                    // LEDs_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> LEDs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                          // LEDs_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> LEDs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                  // LEDs_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> LEDs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [105:0] leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                           // LEDs_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> LEDs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                          // LEDs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> LEDs_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                 // LEDs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> LEDs_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                       // LEDs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> LEDs_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                               // LEDs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> LEDs_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [105:0] leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                        // LEDs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> LEDs_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                       // LEDs_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> LEDs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                     // LEDs_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> LEDs_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                      // LEDs_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> LEDs_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                     // LEDs_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> LEDs_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          switches_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                       // switches_s1_translator:uav_waitrequest -> switches_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] switches_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                        // switches_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> switches_s1_translator:uav_burstcount
	wire   [31:0] switches_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                         // switches_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> switches_s1_translator:uav_writedata
	wire   [31:0] switches_s1_translator_avalon_universal_slave_0_agent_m0_address;                                           // switches_s1_translator_avalon_universal_slave_0_agent:m0_address -> switches_s1_translator:uav_address
	wire          switches_s1_translator_avalon_universal_slave_0_agent_m0_write;                                             // switches_s1_translator_avalon_universal_slave_0_agent:m0_write -> switches_s1_translator:uav_write
	wire          switches_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                              // switches_s1_translator_avalon_universal_slave_0_agent:m0_lock -> switches_s1_translator:uav_lock
	wire          switches_s1_translator_avalon_universal_slave_0_agent_m0_read;                                              // switches_s1_translator_avalon_universal_slave_0_agent:m0_read -> switches_s1_translator:uav_read
	wire   [31:0] switches_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                          // switches_s1_translator:uav_readdata -> switches_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          switches_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                     // switches_s1_translator:uav_readdatavalid -> switches_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          switches_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                       // switches_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> switches_s1_translator:uav_debugaccess
	wire    [3:0] switches_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                        // switches_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> switches_s1_translator:uav_byteenable
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                // switches_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                      // switches_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                              // switches_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [105:0] switches_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                       // switches_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                      // switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> switches_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                             // switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> switches_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                   // switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> switches_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                           // switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> switches_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [105:0] switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                    // switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> switches_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                   // switches_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                 // switches_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> switches_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                  // switches_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> switches_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                 // switches_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> switches_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // jtag_uart_0_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_0_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                       // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_0_avalon_jtag_slave_translator:uav_writedata
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                         // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_0_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                           // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_0_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                            // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_0_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                            // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_0_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                        // jtag_uart_0_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // jtag_uart_0_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_0_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_0_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [105:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [105:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                  // character_lcd_0_avalon_lcd_slave_translator:uav_waitrequest -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                   // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> character_lcd_0_avalon_lcd_slave_translator:uav_burstcount
	wire    [7:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                    // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> character_lcd_0_avalon_lcd_slave_translator:uav_writedata
	wire   [31:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_address;                      // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_address -> character_lcd_0_avalon_lcd_slave_translator:uav_address
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_write;                        // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_write -> character_lcd_0_avalon_lcd_slave_translator:uav_write
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_lock;                         // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_lock -> character_lcd_0_avalon_lcd_slave_translator:uav_lock
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_read;                         // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_read -> character_lcd_0_avalon_lcd_slave_translator:uav_read
	wire    [7:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                     // character_lcd_0_avalon_lcd_slave_translator:uav_readdata -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                // character_lcd_0_avalon_lcd_slave_translator:uav_readdatavalid -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                  // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> character_lcd_0_avalon_lcd_slave_translator:uav_debugaccess
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                   // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> character_lcd_0_avalon_lcd_slave_translator:uav_byteenable
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;           // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                 // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;         // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [78:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                  // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                 // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;        // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;              // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;      // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [78:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;               // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;              // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;            // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire    [7:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;             // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;            // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                    // pixel_buffer_avalon_sram_slave_translator:uav_waitrequest -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                     // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> pixel_buffer_avalon_sram_slave_translator:uav_burstcount
	wire   [15:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                      // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> pixel_buffer_avalon_sram_slave_translator:uav_writedata
	wire   [31:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address;                        // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_address -> pixel_buffer_avalon_sram_slave_translator:uav_address
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write;                          // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_write -> pixel_buffer_avalon_sram_slave_translator:uav_write
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock;                           // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_lock -> pixel_buffer_avalon_sram_slave_translator:uav_lock
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read;                           // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_read -> pixel_buffer_avalon_sram_slave_translator:uav_read
	wire   [15:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                       // pixel_buffer_avalon_sram_slave_translator:uav_readdata -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                  // pixel_buffer_avalon_sram_slave_translator:uav_readdatavalid -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                    // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pixel_buffer_avalon_sram_slave_translator:uav_debugaccess
	wire    [1:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                     // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> pixel_buffer_avalon_sram_slave_translator:uav_byteenable
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;             // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                   // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;           // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [87:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                    // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                   // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;          // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;        // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [87:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                 // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;              // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [15:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;               // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;              // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // pixel_buffer_dma_avalon_control_slave_translator:uav_waitrequest -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> pixel_buffer_dma_avalon_control_slave_translator:uav_burstcount
	wire   [31:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> pixel_buffer_dma_avalon_control_slave_translator:uav_writedata
	wire   [31:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> pixel_buffer_dma_avalon_control_slave_translator:uav_address
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> pixel_buffer_dma_avalon_control_slave_translator:uav_write
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> pixel_buffer_dma_avalon_control_slave_translator:uav_lock
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> pixel_buffer_dma_avalon_control_slave_translator:uav_read
	wire   [31:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // pixel_buffer_dma_avalon_control_slave_translator:uav_readdata -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // pixel_buffer_dma_avalon_control_slave_translator:uav_readdatavalid -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pixel_buffer_dma_avalon_control_slave_translator:uav_debugaccess
	wire    [3:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> pixel_buffer_dma_avalon_control_slave_translator:uav_byteenable
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [105:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [105:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // char_drawer_avalon_char_control_slave_translator:uav_waitrequest -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> char_drawer_avalon_char_control_slave_translator:uav_burstcount
	wire   [31:0] char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> char_drawer_avalon_char_control_slave_translator:uav_writedata
	wire   [31:0] char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> char_drawer_avalon_char_control_slave_translator:uav_address
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> char_drawer_avalon_char_control_slave_translator:uav_write
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> char_drawer_avalon_char_control_slave_translator:uav_lock
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> char_drawer_avalon_char_control_slave_translator:uav_read
	wire   [31:0] char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // char_drawer_avalon_char_control_slave_translator:uav_readdata -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // char_drawer_avalon_char_control_slave_translator:uav_readdatavalid -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> char_drawer_avalon_char_control_slave_translator:uav_debugaccess
	wire    [3:0] char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> char_drawer_avalon_char_control_slave_translator:uav_byteenable
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [105:0] char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [105:0] char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // char_drawer_avalon_char_buffer_slave_translator:uav_waitrequest -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;               // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> char_drawer_avalon_char_buffer_slave_translator:uav_burstcount
	wire    [7:0] char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> char_drawer_avalon_char_buffer_slave_translator:uav_writedata
	wire   [31:0] char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_address;                  // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_address -> char_drawer_avalon_char_buffer_slave_translator:uav_address
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_write;                    // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_write -> char_drawer_avalon_char_buffer_slave_translator:uav_write
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_lock;                     // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_lock -> char_drawer_avalon_char_buffer_slave_translator:uav_lock
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_read;                     // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_read -> char_drawer_avalon_char_buffer_slave_translator:uav_read
	wire    [7:0] char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                 // char_drawer_avalon_char_buffer_slave_translator:uav_readdata -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // char_drawer_avalon_char_buffer_slave_translator:uav_readdatavalid -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> char_drawer_avalon_char_buffer_slave_translator:uav_debugaccess
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;               // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> char_drawer_avalon_char_buffer_slave_translator:uav_byteenable
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;             // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [78:0] char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_data;              // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;             // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [78:0] char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire    [7:0] char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;               // nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                     // nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;             // nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [104:0] nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                      // nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                     // addr_router:sink_ready -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                      // nios2_processor_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_valid;                            // nios2_processor_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                    // nios2_processor_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [104:0] nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_data;                             // nios2_processor_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_ready;                            // addr_router_001:sink_ready -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket;         // pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire          pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_valid;               // pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire          pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket;       // pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire   [86:0] pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_data;                // pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire          pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_ready;               // addr_router_002:sink_ready -> pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                 // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                       // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;               // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [104:0] nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                        // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                       // id_router:sink_ready -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                     // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [104:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                      // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_001:sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                          // sdram_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                // sdram_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                        // sdram_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire   [86:0] sdram_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                 // sdram_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                // id_router_002:sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                           // LEDs_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                 // LEDs_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                         // LEDs_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [104:0] leds_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                  // LEDs_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          leds_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                 // id_router_003:sink_ready -> LEDs_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                       // switches_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                             // switches_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                     // switches_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [104:0] switches_s1_translator_avalon_universal_slave_0_agent_rp_data;                                              // switches_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire          switches_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                             // id_router_004:sink_ready -> switches_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                           // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [104:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                            // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_005:sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                  // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_valid;                        // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire   [77:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_data;                         // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_ready;                        // id_router_006:sink_ready -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                    // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid;                          // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                  // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire   [86:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data;                           // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire          pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready;                          // id_router_007:sink_ready -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [104:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire          pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_008:sink_ready -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire  [104:0] char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire          char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_009:sink_ready -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_valid;                    // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire   [77:0] char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_data;                     // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire          char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_010:sink_ready -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          addr_router_src_endofpacket;                                                                                // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire          addr_router_src_valid;                                                                                      // addr_router:src_valid -> limiter:cmd_sink_valid
	wire          addr_router_src_startofpacket;                                                                              // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [104:0] addr_router_src_data;                                                                                       // addr_router:src_data -> limiter:cmd_sink_data
	wire   [10:0] addr_router_src_channel;                                                                                    // addr_router:src_channel -> limiter:cmd_sink_channel
	wire          addr_router_src_ready;                                                                                      // limiter:cmd_sink_ready -> addr_router:src_ready
	wire          limiter_rsp_src_endofpacket;                                                                                // limiter:rsp_src_endofpacket -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_rsp_src_valid;                                                                                      // limiter:rsp_src_valid -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_rsp_src_startofpacket;                                                                              // limiter:rsp_src_startofpacket -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [104:0] limiter_rsp_src_data;                                                                                       // limiter:rsp_src_data -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [10:0] limiter_rsp_src_channel;                                                                                    // limiter:rsp_src_channel -> nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_rsp_src_ready;                                                                                      // nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire          burst_adapter_source0_endofpacket;                                                                          // burst_adapter:source0_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_source0_valid;                                                                                // burst_adapter:source0_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_source0_startofpacket;                                                                        // burst_adapter:source0_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [86:0] burst_adapter_source0_data;                                                                                 // burst_adapter:source0_data -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_source0_ready;                                                                                // sdram_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire   [10:0] burst_adapter_source0_channel;                                                                              // burst_adapter:source0_channel -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_001_source0_endofpacket;                                                                      // burst_adapter_001:source0_endofpacket -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_001_source0_valid;                                                                            // burst_adapter_001:source0_valid -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_001_source0_startofpacket;                                                                    // burst_adapter_001:source0_startofpacket -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [77:0] burst_adapter_001_source0_data;                                                                             // burst_adapter_001:source0_data -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_001_source0_ready;                                                                            // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	wire   [10:0] burst_adapter_001_source0_channel;                                                                          // burst_adapter_001:source0_channel -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_002_source0_endofpacket;                                                                      // burst_adapter_002:source0_endofpacket -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_002_source0_valid;                                                                            // burst_adapter_002:source0_valid -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_002_source0_startofpacket;                                                                    // burst_adapter_002:source0_startofpacket -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [86:0] burst_adapter_002_source0_data;                                                                             // burst_adapter_002:source0_data -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_002_source0_ready;                                                                            // pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_002:source0_ready
	wire   [10:0] burst_adapter_002_source0_channel;                                                                          // burst_adapter_002:source0_channel -> pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_003_source0_endofpacket;                                                                      // burst_adapter_003:source0_endofpacket -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_003_source0_valid;                                                                            // burst_adapter_003:source0_valid -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_003_source0_startofpacket;                                                                    // burst_adapter_003:source0_startofpacket -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [77:0] burst_adapter_003_source0_data;                                                                             // burst_adapter_003:source0_data -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_003_source0_ready;                                                                            // char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_003:source0_ready
	wire   [10:0] burst_adapter_003_source0_channel;                                                                          // burst_adapter_003:source0_channel -> char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rst_controller_reset_out_reset;                                                                             // rst_controller:reset_out -> [LEDs:reset_n, LEDs_s1_translator:reset, LEDs_s1_translator_avalon_universal_slave_0_agent:reset, LEDs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, addr_router_001:reset, addr_router_002:reset, alpha_blender:reset, burst_adapter:reset, burst_adapter_001:reset, burst_adapter_002:reset, burst_adapter_003:reset, char_drawer:reset, char_drawer_avalon_char_buffer_slave_translator:reset, char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent:reset, char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, char_drawer_avalon_char_control_slave_translator:reset, char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:reset, char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, character_lcd_0:reset, character_lcd_0_avalon_lcd_slave_translator:reset, character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:reset, character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_demux_002:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, cmd_xbar_mux_007:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, irq_mapper:reset, jtag_uart_0:rst_n, jtag_uart_0_avalon_jtag_slave_translator:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter:reset, nios2_processor:reset_n, nios2_processor_data_master_translator:reset, nios2_processor_data_master_translator_avalon_universal_master_0_agent:reset, nios2_processor_instruction_master_translator:reset, nios2_processor_instruction_master_translator_avalon_universal_master_0_agent:reset, nios2_processor_jtag_debug_module_translator:reset, nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, onchip_memory2_0:reset, onchip_memory2_0_s1_translator:reset, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:reset, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pixel_buffer:reset, pixel_buffer_avalon_sram_slave_translator:reset, pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:reset, pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pixel_buffer_dma:reset, pixel_buffer_dma_avalon_control_slave_translator:reset, pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:reset, pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pixel_buffer_dma_avalon_pixel_dma_master_translator:reset, pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:reset, rgb_resampler:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, scaler:reset, sdram:reset_n, sdram_s1_translator:reset, sdram_s1_translator_avalon_universal_slave_0_agent:reset, sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, switches:reset_n, switches_s1_translator:reset, switches_s1_translator_avalon_universal_slave_0_agent:reset, switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, video_fifo:reset_stream_in, width_adapter:reset, width_adapter_001:reset, width_adapter_002:reset, width_adapter_003:reset, width_adapter_004:reset, width_adapter_005:reset, width_adapter_006:reset, width_adapter_007:reset, width_adapter_008:reset, width_adapter_009:reset]
	wire          nios2_processor_jtag_debug_module_reset_reset;                                                              // nios2_processor:jtag_debug_module_resetrequest -> [rst_controller:reset_in0, rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	wire          rst_controller_001_reset_out_reset;                                                                         // rst_controller_001:reset_out -> clocks:reset
	wire          rst_controller_002_reset_out_reset;                                                                         // rst_controller_002:reset_out -> [vga_controller:reset, video_fifo:reset_stream_out]
	wire          cmd_xbar_demux_src0_endofpacket;                                                                            // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                                  // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                          // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [104:0] cmd_xbar_demux_src0_data;                                                                                   // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [10:0] cmd_xbar_demux_src0_channel;                                                                                // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire          cmd_xbar_demux_src0_ready;                                                                                  // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire          cmd_xbar_demux_src1_endofpacket;                                                                            // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                                  // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                          // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [104:0] cmd_xbar_demux_src1_data;                                                                                   // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire   [10:0] cmd_xbar_demux_src1_channel;                                                                                // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire          cmd_xbar_demux_src1_ready;                                                                                  // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                                        // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                              // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                                      // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [104:0] cmd_xbar_demux_001_src0_data;                                                                               // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire   [10:0] cmd_xbar_demux_001_src0_channel;                                                                            // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                                              // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire          cmd_xbar_demux_001_src1_endofpacket;                                                                        // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire          cmd_xbar_demux_001_src1_valid;                                                                              // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire          cmd_xbar_demux_001_src1_startofpacket;                                                                      // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [104:0] cmd_xbar_demux_001_src1_data;                                                                               // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire   [10:0] cmd_xbar_demux_001_src1_channel;                                                                            // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire          cmd_xbar_demux_001_src1_ready;                                                                              // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire          cmd_xbar_demux_001_src3_endofpacket;                                                                        // cmd_xbar_demux_001:src3_endofpacket -> LEDs_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src3_valid;                                                                              // cmd_xbar_demux_001:src3_valid -> LEDs_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src3_startofpacket;                                                                      // cmd_xbar_demux_001:src3_startofpacket -> LEDs_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [104:0] cmd_xbar_demux_001_src3_data;                                                                               // cmd_xbar_demux_001:src3_data -> LEDs_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] cmd_xbar_demux_001_src3_channel;                                                                            // cmd_xbar_demux_001:src3_channel -> LEDs_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src4_endofpacket;                                                                        // cmd_xbar_demux_001:src4_endofpacket -> switches_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src4_valid;                                                                              // cmd_xbar_demux_001:src4_valid -> switches_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src4_startofpacket;                                                                      // cmd_xbar_demux_001:src4_startofpacket -> switches_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [104:0] cmd_xbar_demux_001_src4_data;                                                                               // cmd_xbar_demux_001:src4_data -> switches_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] cmd_xbar_demux_001_src4_channel;                                                                            // cmd_xbar_demux_001:src4_channel -> switches_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src5_endofpacket;                                                                        // cmd_xbar_demux_001:src5_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src5_valid;                                                                              // cmd_xbar_demux_001:src5_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src5_startofpacket;                                                                      // cmd_xbar_demux_001:src5_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [104:0] cmd_xbar_demux_001_src5_data;                                                                               // cmd_xbar_demux_001:src5_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] cmd_xbar_demux_001_src5_channel;                                                                            // cmd_xbar_demux_001:src5_channel -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src8_endofpacket;                                                                        // cmd_xbar_demux_001:src8_endofpacket -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src8_valid;                                                                              // cmd_xbar_demux_001:src8_valid -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src8_startofpacket;                                                                      // cmd_xbar_demux_001:src8_startofpacket -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [104:0] cmd_xbar_demux_001_src8_data;                                                                               // cmd_xbar_demux_001:src8_data -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] cmd_xbar_demux_001_src8_channel;                                                                            // cmd_xbar_demux_001:src8_channel -> pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src9_endofpacket;                                                                        // cmd_xbar_demux_001:src9_endofpacket -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src9_valid;                                                                              // cmd_xbar_demux_001:src9_valid -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src9_startofpacket;                                                                      // cmd_xbar_demux_001:src9_startofpacket -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [104:0] cmd_xbar_demux_001_src9_data;                                                                               // cmd_xbar_demux_001:src9_data -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] cmd_xbar_demux_001_src9_channel;                                                                            // cmd_xbar_demux_001:src9_channel -> char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src0_endofpacket;                                                                        // cmd_xbar_demux_002:src0_endofpacket -> cmd_xbar_mux_007:sink1_endofpacket
	wire          cmd_xbar_demux_002_src0_valid;                                                                              // cmd_xbar_demux_002:src0_valid -> cmd_xbar_mux_007:sink1_valid
	wire          cmd_xbar_demux_002_src0_startofpacket;                                                                      // cmd_xbar_demux_002:src0_startofpacket -> cmd_xbar_mux_007:sink1_startofpacket
	wire   [86:0] cmd_xbar_demux_002_src0_data;                                                                               // cmd_xbar_demux_002:src0_data -> cmd_xbar_mux_007:sink1_data
	wire   [10:0] cmd_xbar_demux_002_src0_channel;                                                                            // cmd_xbar_demux_002:src0_channel -> cmd_xbar_mux_007:sink1_channel
	wire          cmd_xbar_demux_002_src0_ready;                                                                              // cmd_xbar_mux_007:sink1_ready -> cmd_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_src0_endofpacket;                                                                            // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                                  // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                          // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [104:0] rsp_xbar_demux_src0_data;                                                                                   // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [10:0] rsp_xbar_demux_src0_channel;                                                                                // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                                  // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_src1_endofpacket;                                                                            // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire          rsp_xbar_demux_src1_valid;                                                                                  // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire          rsp_xbar_demux_src1_startofpacket;                                                                          // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [104:0] rsp_xbar_demux_src1_data;                                                                                   // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire   [10:0] rsp_xbar_demux_src1_channel;                                                                                // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire          rsp_xbar_demux_src1_ready;                                                                                  // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                                        // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                              // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                                      // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [104:0] rsp_xbar_demux_001_src0_data;                                                                               // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [10:0] rsp_xbar_demux_001_src0_channel;                                                                            // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                              // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_001_src1_endofpacket;                                                                        // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire          rsp_xbar_demux_001_src1_valid;                                                                              // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire          rsp_xbar_demux_001_src1_startofpacket;                                                                      // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [104:0] rsp_xbar_demux_001_src1_data;                                                                               // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire   [10:0] rsp_xbar_demux_001_src1_channel;                                                                            // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire          rsp_xbar_demux_001_src1_ready;                                                                              // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                                        // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                              // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux_001:sink3_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                                      // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [104:0] rsp_xbar_demux_003_src0_data;                                                                               // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux_001:sink3_data
	wire   [10:0] rsp_xbar_demux_003_src0_channel;                                                                            // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux_001:sink3_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                              // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                                        // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                              // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink4_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                                      // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [104:0] rsp_xbar_demux_004_src0_data;                                                                               // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink4_data
	wire   [10:0] rsp_xbar_demux_004_src0_channel;                                                                            // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink4_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                                              // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire          rsp_xbar_demux_005_src0_endofpacket;                                                                        // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire          rsp_xbar_demux_005_src0_valid;                                                                              // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	wire          rsp_xbar_demux_005_src0_startofpacket;                                                                      // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [104:0] rsp_xbar_demux_005_src0_data;                                                                               // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	wire   [10:0] rsp_xbar_demux_005_src0_channel;                                                                            // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	wire          rsp_xbar_demux_005_src0_ready;                                                                              // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire          rsp_xbar_demux_007_src1_endofpacket;                                                                        // rsp_xbar_demux_007:src1_endofpacket -> pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_007_src1_valid;                                                                              // rsp_xbar_demux_007:src1_valid -> pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_007_src1_startofpacket;                                                                      // rsp_xbar_demux_007:src1_startofpacket -> pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [86:0] rsp_xbar_demux_007_src1_data;                                                                               // rsp_xbar_demux_007:src1_data -> pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [10:0] rsp_xbar_demux_007_src1_channel;                                                                            // rsp_xbar_demux_007:src1_channel -> pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_008_src0_endofpacket;                                                                        // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	wire          rsp_xbar_demux_008_src0_valid;                                                                              // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink8_valid
	wire          rsp_xbar_demux_008_src0_startofpacket;                                                                      // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	wire  [104:0] rsp_xbar_demux_008_src0_data;                                                                               // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink8_data
	wire   [10:0] rsp_xbar_demux_008_src0_channel;                                                                            // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink8_channel
	wire          rsp_xbar_demux_008_src0_ready;                                                                              // rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire          rsp_xbar_demux_009_src0_endofpacket;                                                                        // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	wire          rsp_xbar_demux_009_src0_valid;                                                                              // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_001:sink9_valid
	wire          rsp_xbar_demux_009_src0_startofpacket;                                                                      // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	wire  [104:0] rsp_xbar_demux_009_src0_data;                                                                               // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_001:sink9_data
	wire   [10:0] rsp_xbar_demux_009_src0_channel;                                                                            // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_001:sink9_channel
	wire          rsp_xbar_demux_009_src0_ready;                                                                              // rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src0_ready
	wire          limiter_cmd_src_endofpacket;                                                                                // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          limiter_cmd_src_startofpacket;                                                                              // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [104:0] limiter_cmd_src_data;                                                                                       // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire   [10:0] limiter_cmd_src_channel;                                                                                    // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire          limiter_cmd_src_ready;                                                                                      // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                               // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                                     // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                             // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [104:0] rsp_xbar_mux_src_data;                                                                                      // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire   [10:0] rsp_xbar_mux_src_channel;                                                                                   // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire          rsp_xbar_mux_src_ready;                                                                                     // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire          addr_router_001_src_endofpacket;                                                                            // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          addr_router_001_src_valid;                                                                                  // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire          addr_router_001_src_startofpacket;                                                                          // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [104:0] addr_router_001_src_data;                                                                                   // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire   [10:0] addr_router_001_src_channel;                                                                                // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire          addr_router_001_src_ready;                                                                                  // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire          rsp_xbar_mux_001_src_endofpacket;                                                                           // rsp_xbar_mux_001:src_endofpacket -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_001_src_valid;                                                                                 // rsp_xbar_mux_001:src_valid -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_001_src_startofpacket;                                                                         // rsp_xbar_mux_001:src_startofpacket -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [104:0] rsp_xbar_mux_001_src_data;                                                                                  // rsp_xbar_mux_001:src_data -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [10:0] rsp_xbar_mux_001_src_channel;                                                                               // rsp_xbar_mux_001:src_channel -> nios2_processor_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_001_src_ready;                                                                                 // nios2_processor_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	wire          addr_router_002_src_endofpacket;                                                                            // addr_router_002:src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire          addr_router_002_src_valid;                                                                                  // addr_router_002:src_valid -> cmd_xbar_demux_002:sink_valid
	wire          addr_router_002_src_startofpacket;                                                                          // addr_router_002:src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire   [86:0] addr_router_002_src_data;                                                                                   // addr_router_002:src_data -> cmd_xbar_demux_002:sink_data
	wire   [10:0] addr_router_002_src_channel;                                                                                // addr_router_002:src_channel -> cmd_xbar_demux_002:sink_channel
	wire          addr_router_002_src_ready;                                                                                  // cmd_xbar_demux_002:sink_ready -> addr_router_002:src_ready
	wire          rsp_xbar_demux_007_src1_ready;                                                                              // pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_007:src1_ready
	wire          cmd_xbar_mux_src_endofpacket;                                                                               // cmd_xbar_mux:src_endofpacket -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_src_valid;                                                                                     // cmd_xbar_mux:src_valid -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_src_startofpacket;                                                                             // cmd_xbar_mux:src_startofpacket -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [104:0] cmd_xbar_mux_src_data;                                                                                      // cmd_xbar_mux:src_data -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] cmd_xbar_mux_src_channel;                                                                                   // cmd_xbar_mux:src_channel -> nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_src_ready;                                                                                     // nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire          id_router_src_endofpacket;                                                                                  // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                                        // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                                                // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [104:0] id_router_src_data;                                                                                         // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [10:0] id_router_src_channel;                                                                                      // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                                        // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          cmd_xbar_mux_001_src_endofpacket;                                                                           // cmd_xbar_mux_001:src_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_001_src_valid;                                                                                 // cmd_xbar_mux_001:src_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_001_src_startofpacket;                                                                         // cmd_xbar_mux_001:src_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [104:0] cmd_xbar_mux_001_src_data;                                                                                  // cmd_xbar_mux_001:src_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] cmd_xbar_mux_001_src_channel;                                                                               // cmd_xbar_mux_001:src_channel -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_001_src_ready;                                                                                 // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire          id_router_001_src_endofpacket;                                                                              // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          id_router_001_src_valid;                                                                                    // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire          id_router_001_src_startofpacket;                                                                            // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [104:0] id_router_001_src_data;                                                                                     // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire   [10:0] id_router_001_src_channel;                                                                                  // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire          id_router_001_src_ready;                                                                                    // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire          cmd_xbar_mux_002_src_endofpacket;                                                                           // cmd_xbar_mux_002:src_endofpacket -> burst_adapter:sink0_endofpacket
	wire          cmd_xbar_mux_002_src_valid;                                                                                 // cmd_xbar_mux_002:src_valid -> burst_adapter:sink0_valid
	wire          cmd_xbar_mux_002_src_startofpacket;                                                                         // cmd_xbar_mux_002:src_startofpacket -> burst_adapter:sink0_startofpacket
	wire   [86:0] cmd_xbar_mux_002_src_data;                                                                                  // cmd_xbar_mux_002:src_data -> burst_adapter:sink0_data
	wire   [10:0] cmd_xbar_mux_002_src_channel;                                                                               // cmd_xbar_mux_002:src_channel -> burst_adapter:sink0_channel
	wire          cmd_xbar_mux_002_src_ready;                                                                                 // burst_adapter:sink0_ready -> cmd_xbar_mux_002:src_ready
	wire          id_router_002_src_endofpacket;                                                                              // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          id_router_002_src_valid;                                                                                    // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire          id_router_002_src_startofpacket;                                                                            // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire   [86:0] id_router_002_src_data;                                                                                     // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire   [10:0] id_router_002_src_channel;                                                                                  // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire          id_router_002_src_ready;                                                                                    // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire          cmd_xbar_demux_001_src3_ready;                                                                              // LEDs_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src3_ready
	wire          id_router_003_src_endofpacket;                                                                              // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                                    // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                                            // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [104:0] id_router_003_src_data;                                                                                     // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire   [10:0] id_router_003_src_channel;                                                                                  // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                                    // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire          cmd_xbar_demux_001_src4_ready;                                                                              // switches_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src4_ready
	wire          id_router_004_src_endofpacket;                                                                              // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          id_router_004_src_valid;                                                                                    // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire          id_router_004_src_startofpacket;                                                                            // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [104:0] id_router_004_src_data;                                                                                     // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire   [10:0] id_router_004_src_channel;                                                                                  // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire          id_router_004_src_ready;                                                                                    // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire          cmd_xbar_demux_001_src5_ready;                                                                              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src5_ready
	wire          id_router_005_src_endofpacket;                                                                              // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire          id_router_005_src_valid;                                                                                    // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire          id_router_005_src_startofpacket;                                                                            // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [104:0] id_router_005_src_data;                                                                                     // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [10:0] id_router_005_src_channel;                                                                                  // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire          id_router_005_src_ready;                                                                                    // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire          width_adapter_002_src_ready;                                                                                // burst_adapter_001:sink0_ready -> width_adapter_002:out_ready
	wire          id_router_006_src_endofpacket;                                                                              // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire          id_router_006_src_valid;                                                                                    // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire          id_router_006_src_startofpacket;                                                                            // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire   [77:0] id_router_006_src_data;                                                                                     // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire   [10:0] id_router_006_src_channel;                                                                                  // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire          id_router_006_src_ready;                                                                                    // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire          cmd_xbar_mux_007_src_endofpacket;                                                                           // cmd_xbar_mux_007:src_endofpacket -> burst_adapter_002:sink0_endofpacket
	wire          cmd_xbar_mux_007_src_valid;                                                                                 // cmd_xbar_mux_007:src_valid -> burst_adapter_002:sink0_valid
	wire          cmd_xbar_mux_007_src_startofpacket;                                                                         // cmd_xbar_mux_007:src_startofpacket -> burst_adapter_002:sink0_startofpacket
	wire   [86:0] cmd_xbar_mux_007_src_data;                                                                                  // cmd_xbar_mux_007:src_data -> burst_adapter_002:sink0_data
	wire   [10:0] cmd_xbar_mux_007_src_channel;                                                                               // cmd_xbar_mux_007:src_channel -> burst_adapter_002:sink0_channel
	wire          cmd_xbar_mux_007_src_ready;                                                                                 // burst_adapter_002:sink0_ready -> cmd_xbar_mux_007:src_ready
	wire          id_router_007_src_endofpacket;                                                                              // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire          id_router_007_src_valid;                                                                                    // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire          id_router_007_src_startofpacket;                                                                            // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire   [86:0] id_router_007_src_data;                                                                                     // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire   [10:0] id_router_007_src_channel;                                                                                  // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire          id_router_007_src_ready;                                                                                    // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire          cmd_xbar_demux_001_src8_ready;                                                                              // pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src8_ready
	wire          id_router_008_src_endofpacket;                                                                              // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire          id_router_008_src_valid;                                                                                    // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire          id_router_008_src_startofpacket;                                                                            // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [104:0] id_router_008_src_data;                                                                                     // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire   [10:0] id_router_008_src_channel;                                                                                  // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire          id_router_008_src_ready;                                                                                    // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire          cmd_xbar_demux_001_src9_ready;                                                                              // char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src9_ready
	wire          id_router_009_src_endofpacket;                                                                              // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire          id_router_009_src_valid;                                                                                    // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire          id_router_009_src_startofpacket;                                                                            // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [104:0] id_router_009_src_data;                                                                                     // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire   [10:0] id_router_009_src_channel;                                                                                  // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire          id_router_009_src_ready;                                                                                    // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire          width_adapter_004_src_ready;                                                                                // burst_adapter_003:sink0_ready -> width_adapter_004:out_ready
	wire          id_router_010_src_endofpacket;                                                                              // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire          id_router_010_src_valid;                                                                                    // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire          id_router_010_src_startofpacket;                                                                            // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire   [77:0] id_router_010_src_data;                                                                                     // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire   [10:0] id_router_010_src_channel;                                                                                  // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire          id_router_010_src_ready;                                                                                    // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire          cmd_xbar_demux_src2_endofpacket;                                                                            // cmd_xbar_demux:src2_endofpacket -> width_adapter:in_endofpacket
	wire          cmd_xbar_demux_src2_valid;                                                                                  // cmd_xbar_demux:src2_valid -> width_adapter:in_valid
	wire          cmd_xbar_demux_src2_startofpacket;                                                                          // cmd_xbar_demux:src2_startofpacket -> width_adapter:in_startofpacket
	wire  [104:0] cmd_xbar_demux_src2_data;                                                                                   // cmd_xbar_demux:src2_data -> width_adapter:in_data
	wire   [10:0] cmd_xbar_demux_src2_channel;                                                                                // cmd_xbar_demux:src2_channel -> width_adapter:in_channel
	wire          cmd_xbar_demux_src2_ready;                                                                                  // width_adapter:in_ready -> cmd_xbar_demux:src2_ready
	wire          width_adapter_src_endofpacket;                                                                              // width_adapter:out_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire          width_adapter_src_valid;                                                                                    // width_adapter:out_valid -> cmd_xbar_mux_002:sink0_valid
	wire          width_adapter_src_startofpacket;                                                                            // width_adapter:out_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire   [86:0] width_adapter_src_data;                                                                                     // width_adapter:out_data -> cmd_xbar_mux_002:sink0_data
	wire          width_adapter_src_ready;                                                                                    // cmd_xbar_mux_002:sink0_ready -> width_adapter:out_ready
	wire   [10:0] width_adapter_src_channel;                                                                                  // width_adapter:out_channel -> cmd_xbar_mux_002:sink0_channel
	wire          cmd_xbar_demux_001_src2_endofpacket;                                                                        // cmd_xbar_demux_001:src2_endofpacket -> width_adapter_001:in_endofpacket
	wire          cmd_xbar_demux_001_src2_valid;                                                                              // cmd_xbar_demux_001:src2_valid -> width_adapter_001:in_valid
	wire          cmd_xbar_demux_001_src2_startofpacket;                                                                      // cmd_xbar_demux_001:src2_startofpacket -> width_adapter_001:in_startofpacket
	wire  [104:0] cmd_xbar_demux_001_src2_data;                                                                               // cmd_xbar_demux_001:src2_data -> width_adapter_001:in_data
	wire   [10:0] cmd_xbar_demux_001_src2_channel;                                                                            // cmd_xbar_demux_001:src2_channel -> width_adapter_001:in_channel
	wire          cmd_xbar_demux_001_src2_ready;                                                                              // width_adapter_001:in_ready -> cmd_xbar_demux_001:src2_ready
	wire          width_adapter_001_src_endofpacket;                                                                          // width_adapter_001:out_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire          width_adapter_001_src_valid;                                                                                // width_adapter_001:out_valid -> cmd_xbar_mux_002:sink1_valid
	wire          width_adapter_001_src_startofpacket;                                                                        // width_adapter_001:out_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire   [86:0] width_adapter_001_src_data;                                                                                 // width_adapter_001:out_data -> cmd_xbar_mux_002:sink1_data
	wire          width_adapter_001_src_ready;                                                                                // cmd_xbar_mux_002:sink1_ready -> width_adapter_001:out_ready
	wire   [10:0] width_adapter_001_src_channel;                                                                              // width_adapter_001:out_channel -> cmd_xbar_mux_002:sink1_channel
	wire          cmd_xbar_demux_001_src6_endofpacket;                                                                        // cmd_xbar_demux_001:src6_endofpacket -> width_adapter_002:in_endofpacket
	wire          cmd_xbar_demux_001_src6_valid;                                                                              // cmd_xbar_demux_001:src6_valid -> width_adapter_002:in_valid
	wire          cmd_xbar_demux_001_src6_startofpacket;                                                                      // cmd_xbar_demux_001:src6_startofpacket -> width_adapter_002:in_startofpacket
	wire  [104:0] cmd_xbar_demux_001_src6_data;                                                                               // cmd_xbar_demux_001:src6_data -> width_adapter_002:in_data
	wire   [10:0] cmd_xbar_demux_001_src6_channel;                                                                            // cmd_xbar_demux_001:src6_channel -> width_adapter_002:in_channel
	wire          cmd_xbar_demux_001_src6_ready;                                                                              // width_adapter_002:in_ready -> cmd_xbar_demux_001:src6_ready
	wire          width_adapter_002_src_endofpacket;                                                                          // width_adapter_002:out_endofpacket -> burst_adapter_001:sink0_endofpacket
	wire          width_adapter_002_src_valid;                                                                                // width_adapter_002:out_valid -> burst_adapter_001:sink0_valid
	wire          width_adapter_002_src_startofpacket;                                                                        // width_adapter_002:out_startofpacket -> burst_adapter_001:sink0_startofpacket
	wire   [77:0] width_adapter_002_src_data;                                                                                 // width_adapter_002:out_data -> burst_adapter_001:sink0_data
	wire   [10:0] width_adapter_002_src_channel;                                                                              // width_adapter_002:out_channel -> burst_adapter_001:sink0_channel
	wire          cmd_xbar_demux_001_src7_endofpacket;                                                                        // cmd_xbar_demux_001:src7_endofpacket -> width_adapter_003:in_endofpacket
	wire          cmd_xbar_demux_001_src7_valid;                                                                              // cmd_xbar_demux_001:src7_valid -> width_adapter_003:in_valid
	wire          cmd_xbar_demux_001_src7_startofpacket;                                                                      // cmd_xbar_demux_001:src7_startofpacket -> width_adapter_003:in_startofpacket
	wire  [104:0] cmd_xbar_demux_001_src7_data;                                                                               // cmd_xbar_demux_001:src7_data -> width_adapter_003:in_data
	wire   [10:0] cmd_xbar_demux_001_src7_channel;                                                                            // cmd_xbar_demux_001:src7_channel -> width_adapter_003:in_channel
	wire          cmd_xbar_demux_001_src7_ready;                                                                              // width_adapter_003:in_ready -> cmd_xbar_demux_001:src7_ready
	wire          width_adapter_003_src_endofpacket;                                                                          // width_adapter_003:out_endofpacket -> cmd_xbar_mux_007:sink0_endofpacket
	wire          width_adapter_003_src_valid;                                                                                // width_adapter_003:out_valid -> cmd_xbar_mux_007:sink0_valid
	wire          width_adapter_003_src_startofpacket;                                                                        // width_adapter_003:out_startofpacket -> cmd_xbar_mux_007:sink0_startofpacket
	wire   [86:0] width_adapter_003_src_data;                                                                                 // width_adapter_003:out_data -> cmd_xbar_mux_007:sink0_data
	wire          width_adapter_003_src_ready;                                                                                // cmd_xbar_mux_007:sink0_ready -> width_adapter_003:out_ready
	wire   [10:0] width_adapter_003_src_channel;                                                                              // width_adapter_003:out_channel -> cmd_xbar_mux_007:sink0_channel
	wire          cmd_xbar_demux_001_src10_endofpacket;                                                                       // cmd_xbar_demux_001:src10_endofpacket -> width_adapter_004:in_endofpacket
	wire          cmd_xbar_demux_001_src10_valid;                                                                             // cmd_xbar_demux_001:src10_valid -> width_adapter_004:in_valid
	wire          cmd_xbar_demux_001_src10_startofpacket;                                                                     // cmd_xbar_demux_001:src10_startofpacket -> width_adapter_004:in_startofpacket
	wire  [104:0] cmd_xbar_demux_001_src10_data;                                                                              // cmd_xbar_demux_001:src10_data -> width_adapter_004:in_data
	wire   [10:0] cmd_xbar_demux_001_src10_channel;                                                                           // cmd_xbar_demux_001:src10_channel -> width_adapter_004:in_channel
	wire          cmd_xbar_demux_001_src10_ready;                                                                             // width_adapter_004:in_ready -> cmd_xbar_demux_001:src10_ready
	wire          width_adapter_004_src_endofpacket;                                                                          // width_adapter_004:out_endofpacket -> burst_adapter_003:sink0_endofpacket
	wire          width_adapter_004_src_valid;                                                                                // width_adapter_004:out_valid -> burst_adapter_003:sink0_valid
	wire          width_adapter_004_src_startofpacket;                                                                        // width_adapter_004:out_startofpacket -> burst_adapter_003:sink0_startofpacket
	wire   [77:0] width_adapter_004_src_data;                                                                                 // width_adapter_004:out_data -> burst_adapter_003:sink0_data
	wire   [10:0] width_adapter_004_src_channel;                                                                              // width_adapter_004:out_channel -> burst_adapter_003:sink0_channel
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                                        // rsp_xbar_demux_002:src0_endofpacket -> width_adapter_005:in_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                              // rsp_xbar_demux_002:src0_valid -> width_adapter_005:in_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                                      // rsp_xbar_demux_002:src0_startofpacket -> width_adapter_005:in_startofpacket
	wire   [86:0] rsp_xbar_demux_002_src0_data;                                                                               // rsp_xbar_demux_002:src0_data -> width_adapter_005:in_data
	wire   [10:0] rsp_xbar_demux_002_src0_channel;                                                                            // rsp_xbar_demux_002:src0_channel -> width_adapter_005:in_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                              // width_adapter_005:in_ready -> rsp_xbar_demux_002:src0_ready
	wire          width_adapter_005_src_endofpacket;                                                                          // width_adapter_005:out_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire          width_adapter_005_src_valid;                                                                                // width_adapter_005:out_valid -> rsp_xbar_mux:sink2_valid
	wire          width_adapter_005_src_startofpacket;                                                                        // width_adapter_005:out_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [104:0] width_adapter_005_src_data;                                                                                 // width_adapter_005:out_data -> rsp_xbar_mux:sink2_data
	wire          width_adapter_005_src_ready;                                                                                // rsp_xbar_mux:sink2_ready -> width_adapter_005:out_ready
	wire   [10:0] width_adapter_005_src_channel;                                                                              // width_adapter_005:out_channel -> rsp_xbar_mux:sink2_channel
	wire          rsp_xbar_demux_002_src1_endofpacket;                                                                        // rsp_xbar_demux_002:src1_endofpacket -> width_adapter_006:in_endofpacket
	wire          rsp_xbar_demux_002_src1_valid;                                                                              // rsp_xbar_demux_002:src1_valid -> width_adapter_006:in_valid
	wire          rsp_xbar_demux_002_src1_startofpacket;                                                                      // rsp_xbar_demux_002:src1_startofpacket -> width_adapter_006:in_startofpacket
	wire   [86:0] rsp_xbar_demux_002_src1_data;                                                                               // rsp_xbar_demux_002:src1_data -> width_adapter_006:in_data
	wire   [10:0] rsp_xbar_demux_002_src1_channel;                                                                            // rsp_xbar_demux_002:src1_channel -> width_adapter_006:in_channel
	wire          rsp_xbar_demux_002_src1_ready;                                                                              // width_adapter_006:in_ready -> rsp_xbar_demux_002:src1_ready
	wire          width_adapter_006_src_endofpacket;                                                                          // width_adapter_006:out_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire          width_adapter_006_src_valid;                                                                                // width_adapter_006:out_valid -> rsp_xbar_mux_001:sink2_valid
	wire          width_adapter_006_src_startofpacket;                                                                        // width_adapter_006:out_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [104:0] width_adapter_006_src_data;                                                                                 // width_adapter_006:out_data -> rsp_xbar_mux_001:sink2_data
	wire          width_adapter_006_src_ready;                                                                                // rsp_xbar_mux_001:sink2_ready -> width_adapter_006:out_ready
	wire   [10:0] width_adapter_006_src_channel;                                                                              // width_adapter_006:out_channel -> rsp_xbar_mux_001:sink2_channel
	wire          rsp_xbar_demux_006_src0_endofpacket;                                                                        // rsp_xbar_demux_006:src0_endofpacket -> width_adapter_007:in_endofpacket
	wire          rsp_xbar_demux_006_src0_valid;                                                                              // rsp_xbar_demux_006:src0_valid -> width_adapter_007:in_valid
	wire          rsp_xbar_demux_006_src0_startofpacket;                                                                      // rsp_xbar_demux_006:src0_startofpacket -> width_adapter_007:in_startofpacket
	wire   [77:0] rsp_xbar_demux_006_src0_data;                                                                               // rsp_xbar_demux_006:src0_data -> width_adapter_007:in_data
	wire   [10:0] rsp_xbar_demux_006_src0_channel;                                                                            // rsp_xbar_demux_006:src0_channel -> width_adapter_007:in_channel
	wire          rsp_xbar_demux_006_src0_ready;                                                                              // width_adapter_007:in_ready -> rsp_xbar_demux_006:src0_ready
	wire          width_adapter_007_src_endofpacket;                                                                          // width_adapter_007:out_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire          width_adapter_007_src_valid;                                                                                // width_adapter_007:out_valid -> rsp_xbar_mux_001:sink6_valid
	wire          width_adapter_007_src_startofpacket;                                                                        // width_adapter_007:out_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [104:0] width_adapter_007_src_data;                                                                                 // width_adapter_007:out_data -> rsp_xbar_mux_001:sink6_data
	wire          width_adapter_007_src_ready;                                                                                // rsp_xbar_mux_001:sink6_ready -> width_adapter_007:out_ready
	wire   [10:0] width_adapter_007_src_channel;                                                                              // width_adapter_007:out_channel -> rsp_xbar_mux_001:sink6_channel
	wire          rsp_xbar_demux_007_src0_endofpacket;                                                                        // rsp_xbar_demux_007:src0_endofpacket -> width_adapter_008:in_endofpacket
	wire          rsp_xbar_demux_007_src0_valid;                                                                              // rsp_xbar_demux_007:src0_valid -> width_adapter_008:in_valid
	wire          rsp_xbar_demux_007_src0_startofpacket;                                                                      // rsp_xbar_demux_007:src0_startofpacket -> width_adapter_008:in_startofpacket
	wire   [86:0] rsp_xbar_demux_007_src0_data;                                                                               // rsp_xbar_demux_007:src0_data -> width_adapter_008:in_data
	wire   [10:0] rsp_xbar_demux_007_src0_channel;                                                                            // rsp_xbar_demux_007:src0_channel -> width_adapter_008:in_channel
	wire          rsp_xbar_demux_007_src0_ready;                                                                              // width_adapter_008:in_ready -> rsp_xbar_demux_007:src0_ready
	wire          width_adapter_008_src_endofpacket;                                                                          // width_adapter_008:out_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire          width_adapter_008_src_valid;                                                                                // width_adapter_008:out_valid -> rsp_xbar_mux_001:sink7_valid
	wire          width_adapter_008_src_startofpacket;                                                                        // width_adapter_008:out_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [104:0] width_adapter_008_src_data;                                                                                 // width_adapter_008:out_data -> rsp_xbar_mux_001:sink7_data
	wire          width_adapter_008_src_ready;                                                                                // rsp_xbar_mux_001:sink7_ready -> width_adapter_008:out_ready
	wire   [10:0] width_adapter_008_src_channel;                                                                              // width_adapter_008:out_channel -> rsp_xbar_mux_001:sink7_channel
	wire          rsp_xbar_demux_010_src0_endofpacket;                                                                        // rsp_xbar_demux_010:src0_endofpacket -> width_adapter_009:in_endofpacket
	wire          rsp_xbar_demux_010_src0_valid;                                                                              // rsp_xbar_demux_010:src0_valid -> width_adapter_009:in_valid
	wire          rsp_xbar_demux_010_src0_startofpacket;                                                                      // rsp_xbar_demux_010:src0_startofpacket -> width_adapter_009:in_startofpacket
	wire   [77:0] rsp_xbar_demux_010_src0_data;                                                                               // rsp_xbar_demux_010:src0_data -> width_adapter_009:in_data
	wire   [10:0] rsp_xbar_demux_010_src0_channel;                                                                            // rsp_xbar_demux_010:src0_channel -> width_adapter_009:in_channel
	wire          rsp_xbar_demux_010_src0_ready;                                                                              // width_adapter_009:in_ready -> rsp_xbar_demux_010:src0_ready
	wire          width_adapter_009_src_endofpacket;                                                                          // width_adapter_009:out_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	wire          width_adapter_009_src_valid;                                                                                // width_adapter_009:out_valid -> rsp_xbar_mux_001:sink10_valid
	wire          width_adapter_009_src_startofpacket;                                                                        // width_adapter_009:out_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	wire  [104:0] width_adapter_009_src_data;                                                                                 // width_adapter_009:out_data -> rsp_xbar_mux_001:sink10_data
	wire          width_adapter_009_src_ready;                                                                                // rsp_xbar_mux_001:sink10_ready -> width_adapter_009:out_ready
	wire   [10:0] width_adapter_009_src_channel;                                                                              // width_adapter_009:out_channel -> rsp_xbar_mux_001:sink10_channel
	wire   [10:0] limiter_cmd_valid_data;                                                                                     // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire          irq_mapper_receiver0_irq;                                                                                   // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire   [31:0] nios2_processor_d_irq_irq;                                                                                  // irq_mapper:sender_irq -> nios2_processor:d_irq

	nios_system_nios2_processor nios2_processor (
		.clk                                   (clocks_sys_clk_clk),                                                             //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                                //                   reset_n.reset_n
		.d_address                             (nios2_processor_data_master_address),                                            //               data_master.address
		.d_byteenable                          (nios2_processor_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (nios2_processor_data_master_read),                                               //                          .read
		.d_readdata                            (nios2_processor_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (nios2_processor_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (nios2_processor_data_master_write),                                              //                          .write
		.d_writedata                           (nios2_processor_data_master_writedata),                                          //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_processor_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (nios2_processor_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (nios2_processor_instruction_master_read),                                        //                          .read
		.i_readdata                            (nios2_processor_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (nios2_processor_instruction_master_waitrequest),                                 //                          .waitrequest
		.i_readdatavalid                       (nios2_processor_instruction_master_readdatavalid),                               //                          .readdatavalid
		.d_irq                                 (nios2_processor_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_processor_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                                // custom_instruction_master.readra
	);

	nios_system_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clocks_sys_clk_clk),                                            //   clk1.clk
		.address    (onchip_memory2_0_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (onchip_memory2_0_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset)                                 // reset1.reset
	);

	nios_system_switches switches (
		.clk      (clocks_sys_clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                     //               reset.reset_n
		.address  (switches_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (switches_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (switches_export)                                      // external_connection.export
	);

	nios_system_LEDs leds (
		.clk        (clocks_sys_clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (leds_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~leds_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (leds_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (leds_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (leds_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (leds_export)                                        // external_connection.export
	);

	nios_system_jtag_uart_0 jtag_uart_0 (
		.clk            (clocks_sys_clk_clk),                                                       //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                          //             reset.reset_n
		.av_chipselect  (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                                  //               irq.irq
	);

	nios_system_sdram sdram (
		.clk            (clocks_sys_clk_clk),                                    //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                       // reset.reset_n
		.az_addr        (sdram_s1_translator_avalon_anti_slave_0_address),       //    s1.address
		.az_be_n        (~sdram_s1_translator_avalon_anti_slave_0_byteenable),   //      .byteenable_n
		.az_cs          (sdram_s1_translator_avalon_anti_slave_0_chipselect),    //      .chipselect
		.az_data        (sdram_s1_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.az_rd_n        (~sdram_s1_translator_avalon_anti_slave_0_read),         //      .read_n
		.az_wr_n        (~sdram_s1_translator_avalon_anti_slave_0_write),        //      .write_n
		.za_data        (sdram_s1_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.za_valid       (sdram_s1_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.za_waitrequest (sdram_s1_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                                       //  wire.export
		.zs_ba          (sdram_wire_ba),                                         //      .export
		.zs_cas_n       (sdram_wire_cas_n),                                      //      .export
		.zs_cke         (sdram_wire_cke),                                        //      .export
		.zs_cs_n        (sdram_wire_cs_n),                                       //      .export
		.zs_dq          (sdram_wire_dq),                                         //      .export
		.zs_dqm         (sdram_wire_dqm),                                        //      .export
		.zs_ras_n       (sdram_wire_ras_n),                                      //      .export
		.zs_we_n        (sdram_wire_we_n)                                        //      .export
	);

	nios_system_clocks clocks (
		.CLOCK_50    (clk_clk),                            //       clk_in_primary.clk
		.reset       (rst_controller_001_reset_out_reset), // clk_in_primary_reset.reset
		.sys_clk     (clocks_sys_clk_clk),                 //              sys_clk.clk
		.sys_reset_n (),                                   //        sys_clk_reset.reset_n
		.SDRAM_CLK   (sdram_clk_clk),                      //            sdram_clk.clk
		.VGA_CLK     (clocks_vga_clk_clk)                  //              vga_clk.clk
	);

	nios_system_character_lcd_0 character_lcd_0 (
		.clk         (clocks_sys_clk_clk),                                                          //        clock_reset.clk
		.reset       (rst_controller_reset_out_reset),                                              //  clock_reset_reset.reset
		.address     (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_address),     //   avalon_lcd_slave.address
		.chipselect  (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_chipselect),  //                   .chipselect
		.read        (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_read),        //                   .read
		.write       (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_write),       //                   .write
		.writedata   (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_writedata),   //                   .writedata
		.readdata    (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_readdata),    //                   .readdata
		.waitrequest (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_waitrequest), //                   .waitrequest
		.LCD_DATA    (lcd_data_DATA),                                                               // external_interface.export
		.LCD_ON      (lcd_data_ON),                                                                 //                   .export
		.LCD_BLON    (lcd_data_BLON),                                                               //                   .export
		.LCD_EN      (lcd_data_EN),                                                                 //                   .export
		.LCD_RS      (lcd_data_RS),                                                                 //                   .export
		.LCD_RW      (lcd_data_RW)                                                                  //                   .export
	);

	nios_system_pixel_buffer pixel_buffer (
		.clk           (clocks_sys_clk_clk),                                                          //        clock_reset.clk
		.reset         (rst_controller_reset_out_reset),                                              //  clock_reset_reset.reset
		.SRAM_DQ       (sram_DQ),                                                                     // external_interface.export
		.SRAM_ADDR     (sram_ADDR),                                                                   //                   .export
		.SRAM_LB_N     (sram_LB_N),                                                                   //                   .export
		.SRAM_UB_N     (sram_UB_N),                                                                   //                   .export
		.SRAM_CE_N     (sram_CE_N),                                                                   //                   .export
		.SRAM_OE_N     (sram_OE_N),                                                                   //                   .export
		.SRAM_WE_N     (sram_WE_N),                                                                   //                   .export
		.address       (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_address),       //  avalon_sram_slave.address
		.byteenable    (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable),    //                   .byteenable
		.read          (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_read),          //                   .read
		.write         (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_write),         //                   .write
		.writedata     (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_writedata),     //                   .writedata
		.readdata      (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdata),      //                   .readdata
		.readdatavalid (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid)  //                   .readdatavalid
	);

	nios_system_pixel_buffer_dma pixel_buffer_dma (
		.clk                  (clocks_sys_clk_clk),                                                              //             clock_reset.clk
		.reset                (rst_controller_reset_out_reset),                                                  //       clock_reset_reset.reset
		.master_readdatavalid (pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid),                          // avalon_pixel_dma_master.readdatavalid
		.master_waitrequest   (pixel_buffer_dma_avalon_pixel_dma_master_waitrequest),                            //                        .waitrequest
		.master_address       (pixel_buffer_dma_avalon_pixel_dma_master_address),                                //                        .address
		.master_arbiterlock   (pixel_buffer_dma_avalon_pixel_dma_master_lock),                                   //                        .lock
		.master_read          (pixel_buffer_dma_avalon_pixel_dma_master_read),                                   //                        .read
		.master_readdata      (pixel_buffer_dma_avalon_pixel_dma_master_readdata),                               //                        .readdata
		.slave_address        (pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_address),    //    avalon_control_slave.address
		.slave_byteenable     (pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_byteenable), //                        .byteenable
		.slave_read           (pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_read),       //                        .read
		.slave_write          (pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_write),      //                        .write
		.slave_writedata      (pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_writedata),  //                        .writedata
		.slave_readdata       (pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_readdata),   //                        .readdata
		.stream_ready         (pixel_buffer_dma_avalon_pixel_source_ready),                                      //     avalon_pixel_source.ready
		.stream_startofpacket (pixel_buffer_dma_avalon_pixel_source_startofpacket),                              //                        .startofpacket
		.stream_endofpacket   (pixel_buffer_dma_avalon_pixel_source_endofpacket),                                //                        .endofpacket
		.stream_valid         (pixel_buffer_dma_avalon_pixel_source_valid),                                      //                        .valid
		.stream_data          (pixel_buffer_dma_avalon_pixel_source_data)                                        //                        .data
	);

	nios_system_rgb_resampler rgb_resampler (
		.clk                      (clocks_sys_clk_clk),                                 //       clock_reset.clk
		.reset                    (rst_controller_reset_out_reset),                     // clock_reset_reset.reset
		.stream_in_startofpacket  (pixel_buffer_dma_avalon_pixel_source_startofpacket), //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (pixel_buffer_dma_avalon_pixel_source_endofpacket),   //                  .endofpacket
		.stream_in_valid          (pixel_buffer_dma_avalon_pixel_source_valid),         //                  .valid
		.stream_in_ready          (pixel_buffer_dma_avalon_pixel_source_ready),         //                  .ready
		.stream_in_data           (pixel_buffer_dma_avalon_pixel_source_data),          //                  .data
		.stream_out_ready         (rgb_resampler_avalon_rgb_source_ready),              // avalon_rgb_source.ready
		.stream_out_startofpacket (rgb_resampler_avalon_rgb_source_startofpacket),      //                  .startofpacket
		.stream_out_endofpacket   (rgb_resampler_avalon_rgb_source_endofpacket),        //                  .endofpacket
		.stream_out_valid         (rgb_resampler_avalon_rgb_source_valid),              //                  .valid
		.stream_out_data          (rgb_resampler_avalon_rgb_source_data)                //                  .data
	);

	nios_system_scaler scaler (
		.clk                      (clocks_sys_clk_clk),                            //          clock_reset.clk
		.reset                    (rst_controller_reset_out_reset),                //    clock_reset_reset.reset
		.stream_in_startofpacket  (rgb_resampler_avalon_rgb_source_startofpacket), //   avalon_scaler_sink.startofpacket
		.stream_in_endofpacket    (rgb_resampler_avalon_rgb_source_endofpacket),   //                     .endofpacket
		.stream_in_valid          (rgb_resampler_avalon_rgb_source_valid),         //                     .valid
		.stream_in_ready          (rgb_resampler_avalon_rgb_source_ready),         //                     .ready
		.stream_in_data           (rgb_resampler_avalon_rgb_source_data),          //                     .data
		.stream_out_ready         (scaler_avalon_scaler_source_ready),             // avalon_scaler_source.ready
		.stream_out_startofpacket (scaler_avalon_scaler_source_startofpacket),     //                     .startofpacket
		.stream_out_endofpacket   (scaler_avalon_scaler_source_endofpacket),       //                     .endofpacket
		.stream_out_valid         (scaler_avalon_scaler_source_valid),             //                     .valid
		.stream_out_data          (scaler_avalon_scaler_source_data)               //                     .data
	);

	nios_system_video_fifo video_fifo (
		.clk_stream_in            (clocks_sys_clk_clk),                                //         clock_stream_in.clk
		.reset_stream_in          (rst_controller_reset_out_reset),                    //   clock_stream_in_reset.reset
		.clk_stream_out           (clocks_vga_clk_clk),                                //        clock_stream_out.clk
		.reset_stream_out         (rst_controller_002_reset_out_reset),                //  clock_stream_out_reset.reset
		.stream_in_ready          (alpha_blender_avalon_blended_source_ready),         //   avalon_dc_buffer_sink.ready
		.stream_in_startofpacket  (alpha_blender_avalon_blended_source_startofpacket), //                        .startofpacket
		.stream_in_endofpacket    (alpha_blender_avalon_blended_source_endofpacket),   //                        .endofpacket
		.stream_in_valid          (alpha_blender_avalon_blended_source_valid),         //                        .valid
		.stream_in_data           (alpha_blender_avalon_blended_source_data),          //                        .data
		.stream_out_ready         (video_fifo_avalon_dc_buffer_source_ready),          // avalon_dc_buffer_source.ready
		.stream_out_startofpacket (video_fifo_avalon_dc_buffer_source_startofpacket),  //                        .startofpacket
		.stream_out_endofpacket   (video_fifo_avalon_dc_buffer_source_endofpacket),    //                        .endofpacket
		.stream_out_valid         (video_fifo_avalon_dc_buffer_source_valid),          //                        .valid
		.stream_out_data          (video_fifo_avalon_dc_buffer_source_data)            //                        .data
	);

	nios_system_vga_controller vga_controller (
		.clk           (clocks_vga_clk_clk),                               //        clock_reset.clk
		.reset         (rst_controller_002_reset_out_reset),               //  clock_reset_reset.reset
		.data          (video_fifo_avalon_dc_buffer_source_data),          //    avalon_vga_sink.data
		.startofpacket (video_fifo_avalon_dc_buffer_source_startofpacket), //                   .startofpacket
		.endofpacket   (video_fifo_avalon_dc_buffer_source_endofpacket),   //                   .endofpacket
		.valid         (video_fifo_avalon_dc_buffer_source_valid),         //                   .valid
		.ready         (video_fifo_avalon_dc_buffer_source_ready),         //                   .ready
		.VGA_CLK       (vga_controller_CLK),                               // external_interface.export
		.VGA_HS        (vga_controller_HS),                                //                   .export
		.VGA_VS        (vga_controller_VS),                                //                   .export
		.VGA_BLANK     (vga_controller_BLANK),                             //                   .export
		.VGA_SYNC      (vga_controller_SYNC),                              //                   .export
		.VGA_R         (vga_controller_R),                                 //                   .export
		.VGA_G         (vga_controller_G),                                 //                   .export
		.VGA_B         (vga_controller_B)                                  //                   .export
	);

	nios_system_char_drawer char_drawer (
		.clk                  (clocks_sys_clk_clk),                                                              //               clock_reset.clk
		.reset                (rst_controller_reset_out_reset),                                                  //         clock_reset_reset.reset
		.ctrl_address         (char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_address),    // avalon_char_control_slave.address
		.ctrl_byteenable      (char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_byteenable), //                          .byteenable
		.ctrl_chipselect      (char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_chipselect), //                          .chipselect
		.ctrl_read            (char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_read),       //                          .read
		.ctrl_write           (char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_write),      //                          .write
		.ctrl_writedata       (char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_writedata),  //                          .writedata
		.ctrl_readdata        (char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_readdata),   //                          .readdata
		.buf_byteenable       (char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_byteenable),  //  avalon_char_buffer_slave.byteenable
		.buf_chipselect       (char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_chipselect),  //                          .chipselect
		.buf_read             (char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_read),        //                          .read
		.buf_write            (char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_write),       //                          .write
		.buf_writedata        (char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_writedata),   //                          .writedata
		.buf_readdata         (char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_readdata),    //                          .readdata
		.buf_waitrequest      (char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_waitrequest), //                          .waitrequest
		.buf_address          (char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_address),     //                          .address
		.stream_ready         (char_drawer_avalon_char_source_ready),                                            //        avalon_char_source.ready
		.stream_startofpacket (char_drawer_avalon_char_source_startofpacket),                                    //                          .startofpacket
		.stream_endofpacket   (char_drawer_avalon_char_source_endofpacket),                                      //                          .endofpacket
		.stream_valid         (char_drawer_avalon_char_source_valid),                                            //                          .valid
		.stream_data          (char_drawer_avalon_char_source_data)                                              //                          .data
	);

	nios_system_alpha_blender alpha_blender (
		.clk                      (clocks_sys_clk_clk),                                //            clock_reset.clk
		.reset                    (rst_controller_reset_out_reset),                    //      clock_reset_reset.reset
		.foreground_data          (char_drawer_avalon_char_source_data),               // avalon_foreground_sink.data
		.foreground_startofpacket (char_drawer_avalon_char_source_startofpacket),      //                       .startofpacket
		.foreground_endofpacket   (char_drawer_avalon_char_source_endofpacket),        //                       .endofpacket
		.foreground_valid         (char_drawer_avalon_char_source_valid),              //                       .valid
		.foreground_ready         (char_drawer_avalon_char_source_ready),              //                       .ready
		.background_data          (scaler_avalon_scaler_source_data),                  // avalon_background_sink.data
		.background_startofpacket (scaler_avalon_scaler_source_startofpacket),         //                       .startofpacket
		.background_endofpacket   (scaler_avalon_scaler_source_endofpacket),           //                       .endofpacket
		.background_valid         (scaler_avalon_scaler_source_valid),                 //                       .valid
		.background_ready         (scaler_avalon_scaler_source_ready),                 //                       .ready
		.output_ready             (alpha_blender_avalon_blended_source_ready),         //  avalon_blended_source.ready
		.output_data              (alpha_blender_avalon_blended_source_data),          //                       .data
		.output_startofpacket     (alpha_blender_avalon_blended_source_startofpacket), //                       .startofpacket
		.output_endofpacket       (alpha_blender_avalon_blended_source_endofpacket),   //                       .endofpacket
		.output_valid             (alpha_blender_avalon_blended_source_valid)          //                       .valid
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (25),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_processor_instruction_master_translator (
		.clk                   (clocks_sys_clk_clk),                                                                    //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                        //                     reset.reset
		.uav_address           (nios2_processor_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (nios2_processor_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (nios2_processor_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (nios2_processor_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (nios2_processor_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (nios2_processor_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (nios2_processor_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (nios2_processor_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (nios2_processor_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (nios2_processor_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (nios2_processor_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (nios2_processor_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (nios2_processor_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (nios2_processor_instruction_master_read),                                               //                          .read
		.av_readdata           (nios2_processor_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (nios2_processor_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                                  //               (terminated)
		.av_byteenable         (4'b1111),                                                                               //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                                  //               (terminated)
		.av_begintransfer      (1'b0),                                                                                  //               (terminated)
		.av_chipselect         (1'b0),                                                                                  //               (terminated)
		.av_write              (1'b0),                                                                                  //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                                  //               (terminated)
		.av_lock               (1'b0),                                                                                  //               (terminated)
		.av_debugaccess        (1'b0),                                                                                  //               (terminated)
		.uav_clken             (),                                                                                      //               (terminated)
		.av_clken              (1'b1)                                                                                   //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (25),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_processor_data_master_translator (
		.clk                   (clocks_sys_clk_clk),                                                             //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                 //                     reset.reset
		.uav_address           (nios2_processor_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (nios2_processor_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (nios2_processor_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (nios2_processor_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (nios2_processor_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (nios2_processor_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (nios2_processor_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (nios2_processor_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (nios2_processor_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (nios2_processor_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (nios2_processor_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (nios2_processor_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (nios2_processor_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (nios2_processor_data_master_byteenable),                                         //                          .byteenable
		.av_read               (nios2_processor_data_master_read),                                               //                          .read
		.av_readdata           (nios2_processor_data_master_readdata),                                           //                          .readdata
		.av_write              (nios2_processor_data_master_write),                                              //                          .write
		.av_writedata          (nios2_processor_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (nios2_processor_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                                           //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                           //               (terminated)
		.av_begintransfer      (1'b0),                                                                           //               (terminated)
		.av_chipselect         (1'b0),                                                                           //               (terminated)
		.av_readdatavalid      (),                                                                               //               (terminated)
		.av_lock               (1'b0),                                                                           //               (terminated)
		.uav_clken             (),                                                                               //               (terminated)
		.av_clken              (1'b1)                                                                            //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (16),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (2),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (2),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (2),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) pixel_buffer_dma_avalon_pixel_dma_master_translator (
		.clk                   (clocks_sys_clk_clk),                                                                          //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                              //                     reset.reset
		.uav_address           (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (pixel_buffer_dma_avalon_pixel_dma_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (pixel_buffer_dma_avalon_pixel_dma_master_waitrequest),                                        //                          .waitrequest
		.av_read               (pixel_buffer_dma_avalon_pixel_dma_master_read),                                               //                          .read
		.av_readdata           (pixel_buffer_dma_avalon_pixel_dma_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid),                                      //                          .readdatavalid
		.av_lock               (pixel_buffer_dma_avalon_pixel_dma_master_lock),                                               //                          .lock
		.av_burstcount         (1'b1),                                                                                        //               (terminated)
		.av_byteenable         (2'b11),                                                                                       //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                                        //               (terminated)
		.av_begintransfer      (1'b0),                                                                                        //               (terminated)
		.av_chipselect         (1'b0),                                                                                        //               (terminated)
		.av_write              (1'b0),                                                                                        //               (terminated)
		.av_writedata          (16'b0000000000000000),                                                                        //               (terminated)
		.av_debugaccess        (1'b0),                                                                                        //               (terminated)
		.uav_clken             (),                                                                                            //               (terminated)
		.av_clken              (1'b1)                                                                                         //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) nios2_processor_jtag_debug_module_translator (
		.clk                   (clocks_sys_clk_clk),                                                                           //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                               //                    reset.reset
		.uav_address           (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (nios2_processor_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                                             //              (terminated)
		.av_burstcount         (),                                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                         //              (terminated)
		.av_waitrequest        (1'b0),                                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                                             //              (terminated)
		.av_lock               (),                                                                                             //              (terminated)
		.av_clken              (),                                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                                         //              (terminated)
		.av_outputenable       ()                                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (10),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) onchip_memory2_0_s1_translator (
		.clk                   (clocks_sys_clk_clk),                                                             //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                 //                    reset.reset
		.uav_address           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (onchip_memory2_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (onchip_memory2_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                               //              (terminated)
		.av_begintransfer      (),                                                                               //              (terminated)
		.av_beginbursttransfer (),                                                                               //              (terminated)
		.av_burstcount         (),                                                                               //              (terminated)
		.av_readdatavalid      (1'b0),                                                                           //              (terminated)
		.av_waitrequest        (1'b0),                                                                           //              (terminated)
		.av_writebyteenable    (),                                                                               //              (terminated)
		.av_lock               (),                                                                               //              (terminated)
		.uav_clken             (1'b0),                                                                           //              (terminated)
		.av_debugaccess        (),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (22),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sdram_s1_translator (
		.clk                   (clocks_sys_clk_clk),                                                  //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                      //                    reset.reset
		.uav_address           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sdram_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sdram_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sdram_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sdram_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sdram_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sdram_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (sdram_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (sdram_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (sdram_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (sdram_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                    //              (terminated)
		.av_beginbursttransfer (),                                                                    //              (terminated)
		.av_burstcount         (),                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                    //              (terminated)
		.av_lock               (),                                                                    //              (terminated)
		.av_clken              (),                                                                    //              (terminated)
		.uav_clken             (1'b0),                                                                //              (terminated)
		.av_debugaccess        (),                                                                    //              (terminated)
		.av_outputenable       ()                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) leds_s1_translator (
		.clk                   (clocks_sys_clk_clk),                                                 //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address           (leds_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (leds_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (leds_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (leds_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (leds_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (leds_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (leds_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (leds_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (leds_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                   //              (terminated)
		.av_begintransfer      (),                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                   //              (terminated)
		.av_burstcount         (),                                                                   //              (terminated)
		.av_byteenable         (),                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                               //              (terminated)
		.av_writebyteenable    (),                                                                   //              (terminated)
		.av_lock               (),                                                                   //              (terminated)
		.av_clken              (),                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                               //              (terminated)
		.av_debugaccess        (),                                                                   //              (terminated)
		.av_outputenable       ()                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) switches_s1_translator (
		.clk                   (clocks_sys_clk_clk),                                                     //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                         //                    reset.reset
		.uav_address           (switches_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (switches_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (switches_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (switches_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (switches_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (switches_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (switches_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (switches_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (switches_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (switches_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (switches_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (switches_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata           (switches_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write              (),                                                                       //              (terminated)
		.av_read               (),                                                                       //              (terminated)
		.av_writedata          (),                                                                       //              (terminated)
		.av_begintransfer      (),                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                       //              (terminated)
		.av_burstcount         (),                                                                       //              (terminated)
		.av_byteenable         (),                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                   //              (terminated)
		.av_waitrequest        (1'b0),                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                       //              (terminated)
		.av_lock               (),                                                                       //              (terminated)
		.av_chipselect         (),                                                                       //              (terminated)
		.av_clken              (),                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                   //              (terminated)
		.av_debugaccess        (),                                                                       //              (terminated)
		.av_outputenable       ()                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_0_avalon_jtag_slave_translator (
		.clk                   (clocks_sys_clk_clk),                                                                       //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                           //                    reset.reset
		.uav_address           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                                         //              (terminated)
		.av_burstcount         (),                                                                                         //              (terminated)
		.av_byteenable         (),                                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                                         //              (terminated)
		.av_lock               (),                                                                                         //              (terminated)
		.av_clken              (),                                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                                     //              (terminated)
		.av_debugaccess        (),                                                                                         //              (terminated)
		.av_outputenable       ()                                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) character_lcd_0_avalon_lcd_slave_translator (
		.clk                   (clocks_sys_clk_clk),                                                                          //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                              //                    reset.reset
		.uav_address           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                            //              (terminated)
		.av_beginbursttransfer (),                                                                                            //              (terminated)
		.av_burstcount         (),                                                                                            //              (terminated)
		.av_byteenable         (),                                                                                            //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                        //              (terminated)
		.av_writebyteenable    (),                                                                                            //              (terminated)
		.av_lock               (),                                                                                            //              (terminated)
		.av_clken              (),                                                                                            //              (terminated)
		.uav_clken             (1'b0),                                                                                        //              (terminated)
		.av_debugaccess        (),                                                                                            //              (terminated)
		.av_outputenable       ()                                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (18),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pixel_buffer_avalon_sram_slave_translator (
		.clk                   (clocks_sys_clk_clk),                                                                        //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                            //                    reset.reset
		.uav_address           (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_begintransfer      (),                                                                                          //              (terminated)
		.av_beginbursttransfer (),                                                                                          //              (terminated)
		.av_burstcount         (),                                                                                          //              (terminated)
		.av_waitrequest        (1'b0),                                                                                      //              (terminated)
		.av_writebyteenable    (),                                                                                          //              (terminated)
		.av_lock               (),                                                                                          //              (terminated)
		.av_chipselect         (),                                                                                          //              (terminated)
		.av_clken              (),                                                                                          //              (terminated)
		.uav_clken             (1'b0),                                                                                      //              (terminated)
		.av_debugaccess        (),                                                                                          //              (terminated)
		.av_outputenable       ()                                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pixel_buffer_dma_avalon_control_slave_translator (
		.clk                   (clocks_sys_clk_clk),                                                                               //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                                   //                    reset.reset
		.uav_address           (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_begintransfer      (),                                                                                                 //              (terminated)
		.av_beginbursttransfer (),                                                                                                 //              (terminated)
		.av_burstcount         (),                                                                                                 //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                             //              (terminated)
		.av_waitrequest        (1'b0),                                                                                             //              (terminated)
		.av_writebyteenable    (),                                                                                                 //              (terminated)
		.av_lock               (),                                                                                                 //              (terminated)
		.av_chipselect         (),                                                                                                 //              (terminated)
		.av_clken              (),                                                                                                 //              (terminated)
		.uav_clken             (1'b0),                                                                                             //              (terminated)
		.av_debugaccess        (),                                                                                                 //              (terminated)
		.av_outputenable       ()                                                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) char_drawer_avalon_char_control_slave_translator (
		.clk                   (clocks_sys_clk_clk),                                                                               //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                                   //                    reset.reset
		.uav_address           (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (char_drawer_avalon_char_control_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                                 //              (terminated)
		.av_beginbursttransfer (),                                                                                                 //              (terminated)
		.av_burstcount         (),                                                                                                 //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                             //              (terminated)
		.av_waitrequest        (1'b0),                                                                                             //              (terminated)
		.av_writebyteenable    (),                                                                                                 //              (terminated)
		.av_lock               (),                                                                                                 //              (terminated)
		.av_clken              (),                                                                                                 //              (terminated)
		.uav_clken             (1'b0),                                                                                             //              (terminated)
		.av_debugaccess        (),                                                                                                 //              (terminated)
		.av_outputenable       ()                                                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (13),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) char_drawer_avalon_char_buffer_slave_translator (
		.clk                   (clocks_sys_clk_clk),                                                                              //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                                  //                    reset.reset
		.uav_address           (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (char_drawer_avalon_char_buffer_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                                //              (terminated)
		.av_burstcount         (),                                                                                                //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                            //              (terminated)
		.av_writebyteenable    (),                                                                                                //              (terminated)
		.av_lock               (),                                                                                                //              (terminated)
		.av_clken              (),                                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                                            //              (terminated)
		.av_debugaccess        (),                                                                                                //              (terminated)
		.av_outputenable       ()                                                                                                 //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (98),
		.PKT_PROTECTION_L          (96),
		.PKT_BEGIN_BURST           (86),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (94),
		.PKT_DEST_ID_L             (91),
		.PKT_THREAD_ID_H           (95),
		.PKT_THREAD_ID_L           (95),
		.PKT_CACHE_H               (102),
		.PKT_CACHE_L               (99),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.ST_DATA_W                 (105),
		.ST_CHANNEL_W              (11),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (4'b0000)
	) nios2_processor_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (clocks_sys_clk_clk),                                                                             //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                                 // clk_reset.reset
		.av_address       (nios2_processor_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (nios2_processor_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (nios2_processor_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (nios2_processor_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (nios2_processor_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (nios2_processor_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (nios2_processor_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (nios2_processor_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (nios2_processor_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (nios2_processor_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (nios2_processor_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_rsp_src_valid),                                                                          //        rp.valid
		.rp_data          (limiter_rsp_src_data),                                                                           //          .data
		.rp_channel       (limiter_rsp_src_channel),                                                                        //          .channel
		.rp_startofpacket (limiter_rsp_src_startofpacket),                                                                  //          .startofpacket
		.rp_endofpacket   (limiter_rsp_src_endofpacket),                                                                    //          .endofpacket
		.rp_ready         (limiter_rsp_src_ready)                                                                           //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (98),
		.PKT_PROTECTION_L          (96),
		.PKT_BEGIN_BURST           (86),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (94),
		.PKT_DEST_ID_L             (91),
		.PKT_THREAD_ID_H           (95),
		.PKT_THREAD_ID_L           (95),
		.PKT_CACHE_H               (102),
		.PKT_CACHE_L               (99),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.ST_DATA_W                 (105),
		.ST_CHANNEL_W              (11),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) nios2_processor_data_master_translator_avalon_universal_master_0_agent (
		.clk              (clocks_sys_clk_clk),                                                                      //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.av_address       (nios2_processor_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (nios2_processor_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (nios2_processor_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (nios2_processor_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (nios2_processor_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (nios2_processor_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (nios2_processor_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (nios2_processor_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (nios2_processor_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (nios2_processor_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (nios2_processor_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_001_src_valid),                                                              //        rp.valid
		.rp_data          (rsp_xbar_mux_001_src_data),                                                               //          .data
		.rp_channel       (rsp_xbar_mux_001_src_channel),                                                            //          .channel
		.rp_startofpacket (rsp_xbar_mux_001_src_startofpacket),                                                      //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_001_src_endofpacket),                                                        //          .endofpacket
		.rp_ready         (rsp_xbar_mux_001_src_ready)                                                               //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (80),
		.PKT_PROTECTION_L          (78),
		.PKT_BEGIN_BURST           (68),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_SRC_ID_H              (72),
		.PKT_SRC_ID_L              (69),
		.PKT_DEST_ID_H             (76),
		.PKT_DEST_ID_L             (73),
		.PKT_THREAD_ID_H           (77),
		.PKT_THREAD_ID_L           (77),
		.PKT_CACHE_H               (84),
		.PKT_CACHE_L               (81),
		.PKT_ADDR_SIDEBAND_H       (67),
		.PKT_ADDR_SIDEBAND_L       (67),
		.ST_DATA_W                 (87),
		.ST_CHANNEL_W              (11),
		.AV_BURSTCOUNT_W           (2),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (2),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent (
		.clk              (clocks_sys_clk_clk),                                                                                   //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                                       // clk_reset.reset
		.av_address       (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_demux_007_src1_valid),                                                                        //        rp.valid
		.rp_data          (rsp_xbar_demux_007_src1_data),                                                                         //          .data
		.rp_channel       (rsp_xbar_demux_007_src1_channel),                                                                      //          .channel
		.rp_startofpacket (rsp_xbar_demux_007_src1_startofpacket),                                                                //          .startofpacket
		.rp_endofpacket   (rsp_xbar_demux_007_src1_endofpacket),                                                                  //          .endofpacket
		.rp_ready         (rsp_xbar_demux_007_src1_ready)                                                                         //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (94),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (98),
		.PKT_PROTECTION_L          (96),
		.PKT_RESPONSE_STATUS_H     (104),
		.PKT_RESPONSE_STATUS_L     (103),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (105),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                                     //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                         //       clk_reset.reset
		.m0_address              (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                                 //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                                 //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                                  //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                           //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                               //                .channel
		.rf_sink_ready           (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (106),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                                     //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                         // clk_reset.reset
		.in_data           (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                                   // (terminated)
		.csr_readdata      (),                                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                   // (terminated)
		.almost_full_data  (),                                                                                                       // (terminated)
		.almost_empty_data (),                                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                                   // (terminated)
		.out_empty         (),                                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                                   // (terminated)
		.out_error         (),                                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                                   // (terminated)
		.out_channel       ()                                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (94),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (98),
		.PKT_PROTECTION_L          (96),
		.PKT_RESPONSE_STATUS_H     (104),
		.PKT_RESPONSE_STATUS_L     (103),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (105),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                       //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                               //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                               //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                                //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                                         //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                             //                .channel
		.rf_sink_ready           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (106),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                       //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (68),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (72),
		.PKT_SRC_ID_L              (69),
		.PKT_DEST_ID_H             (76),
		.PKT_DEST_ID_L             (73),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (80),
		.PKT_PROTECTION_L          (78),
		.PKT_RESPONSE_STATUS_H     (86),
		.PKT_RESPONSE_STATUS_L     (85),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (87),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sdram_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                            //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sdram_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sdram_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                   //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                   //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                    //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                             //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                 //                .channel
		.rf_sink_ready           (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (88),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                            //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.in_data           (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (94),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (98),
		.PKT_PROTECTION_L          (96),
		.PKT_RESPONSE_STATUS_H     (104),
		.PKT_RESPONSE_STATUS_L     (103),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (105),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) leds_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (leds_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (leds_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (leds_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (leds_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (leds_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (leds_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (leds_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src3_ready),                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src3_valid),                                                //                .valid
		.cp_data                 (cmd_xbar_demux_001_src3_data),                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src3_startofpacket),                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src3_endofpacket),                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src3_channel),                                              //                .channel
		.rf_sink_ready           (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (106),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (94),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (98),
		.PKT_PROTECTION_L          (96),
		.PKT_RESPONSE_STATUS_H     (104),
		.PKT_RESPONSE_STATUS_L     (103),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (105),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) switches_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                               //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                   //       clk_reset.reset
		.m0_address              (switches_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (switches_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (switches_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (switches_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (switches_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (switches_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (switches_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (switches_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (switches_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (switches_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (switches_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (switches_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (switches_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (switches_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (switches_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (switches_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src4_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src4_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src4_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src4_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src4_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src4_channel),                                                  //                .channel
		.rf_sink_ready           (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (switches_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (106),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.in_data           (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (switches_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (switches_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (94),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (98),
		.PKT_PROTECTION_L          (96),
		.PKT_RESPONSE_STATUS_H     (104),
		.PKT_RESPONSE_STATUS_L     (103),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (105),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                     //       clk_reset.reset
		.m0_address              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src5_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src5_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_001_src5_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src5_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src5_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src5_channel),                                                                    //                .channel
		.rf_sink_ready           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (106),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                     // clk_reset.reset
		.in_data           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (59),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (63),
		.PKT_SRC_ID_L              (60),
		.PKT_DEST_ID_H             (67),
		.PKT_DEST_ID_L             (64),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_PROTECTION_H          (71),
		.PKT_PROTECTION_L          (69),
		.PKT_RESPONSE_STATUS_H     (77),
		.PKT_RESPONSE_STATUS_L     (76),
		.PKT_BURST_SIZE_H          (55),
		.PKT_BURST_SIZE_L          (53),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (78),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                                    //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                        //       clk_reset.reset
		.m0_address              (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_001_source0_ready),                                                                       //              cp.ready
		.cp_valid                (burst_adapter_001_source0_valid),                                                                       //                .valid
		.cp_data                 (burst_adapter_001_source0_data),                                                                        //                .data
		.cp_startofpacket        (burst_adapter_001_source0_startofpacket),                                                               //                .startofpacket
		.cp_endofpacket          (burst_adapter_001_source0_endofpacket),                                                                 //                .endofpacket
		.cp_channel              (burst_adapter_001_source0_channel),                                                                     //                .channel
		.rf_sink_ready           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (79),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                                    //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                        // clk_reset.reset
		.in_data           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                                  // (terminated)
		.csr_readdata      (),                                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                  // (terminated)
		.almost_full_data  (),                                                                                                      // (terminated)
		.almost_empty_data (),                                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                                  // (terminated)
		.out_empty         (),                                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                                  // (terminated)
		.out_error         (),                                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                                  // (terminated)
		.out_channel       ()                                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (68),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (72),
		.PKT_SRC_ID_L              (69),
		.PKT_DEST_ID_H             (76),
		.PKT_DEST_ID_L             (73),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (80),
		.PKT_PROTECTION_L          (78),
		.PKT_RESPONSE_STATUS_H     (86),
		.PKT_RESPONSE_STATUS_L     (85),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (87),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                      //       clk_reset.reset
		.m0_address              (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_002_source0_ready),                                                                     //              cp.ready
		.cp_valid                (burst_adapter_002_source0_valid),                                                                     //                .valid
		.cp_data                 (burst_adapter_002_source0_data),                                                                      //                .data
		.cp_startofpacket        (burst_adapter_002_source0_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (burst_adapter_002_source0_endofpacket),                                                               //                .endofpacket
		.cp_channel              (burst_adapter_002_source0_channel),                                                                   //                .channel
		.rf_sink_ready           (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (88),
		.FIFO_DEPTH          (3),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                      // clk_reset.reset
		.in_data           (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                                // (terminated)
		.csr_readdata      (),                                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                // (terminated)
		.almost_full_data  (),                                                                                                    // (terminated)
		.almost_empty_data (),                                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                                // (terminated)
		.out_empty         (),                                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                                // (terminated)
		.out_error         (),                                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                                // (terminated)
		.out_channel       ()                                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (94),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (98),
		.PKT_PROTECTION_L          (96),
		.PKT_RESPONSE_STATUS_H     (104),
		.PKT_RESPONSE_STATUS_L     (103),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (105),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                                         //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                             //       clk_reset.reset
		.m0_address              (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src8_ready),                                                                              //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src8_valid),                                                                              //                .valid
		.cp_data                 (cmd_xbar_demux_001_src8_data),                                                                               //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src8_startofpacket),                                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src8_endofpacket),                                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src8_channel),                                                                            //                .channel
		.rf_sink_ready           (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (106),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                                         //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                             // clk_reset.reset
		.in_data           (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                                       // (terminated)
		.csr_readdata      (),                                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                       // (terminated)
		.almost_full_data  (),                                                                                                           // (terminated)
		.almost_empty_data (),                                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                                       // (terminated)
		.out_empty         (),                                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                                       // (terminated)
		.out_error         (),                                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                                       // (terminated)
		.out_channel       ()                                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (94),
		.PKT_DEST_ID_L             (91),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (98),
		.PKT_PROTECTION_L          (96),
		.PKT_RESPONSE_STATUS_H     (104),
		.PKT_RESPONSE_STATUS_L     (103),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (105),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                                         //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                             //       clk_reset.reset
		.m0_address              (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src9_ready),                                                                              //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src9_valid),                                                                              //                .valid
		.cp_data                 (cmd_xbar_demux_001_src9_data),                                                                               //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src9_startofpacket),                                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src9_endofpacket),                                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src9_channel),                                                                            //                .channel
		.rf_sink_ready           (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (106),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                                         //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                             // clk_reset.reset
		.in_data           (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                                       // (terminated)
		.csr_readdata      (),                                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                       // (terminated)
		.almost_full_data  (),                                                                                                           // (terminated)
		.almost_empty_data (),                                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                                       // (terminated)
		.out_empty         (),                                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                                       // (terminated)
		.out_error         (),                                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                                       // (terminated)
		.out_channel       ()                                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (59),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (63),
		.PKT_SRC_ID_L              (60),
		.PKT_DEST_ID_H             (67),
		.PKT_DEST_ID_L             (64),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_PROTECTION_H          (71),
		.PKT_PROTECTION_L          (69),
		.PKT_RESPONSE_STATUS_H     (77),
		.PKT_RESPONSE_STATUS_L     (76),
		.PKT_BURST_SIZE_H          (55),
		.PKT_BURST_SIZE_L          (53),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (78),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clocks_sys_clk_clk),                                                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                            //       clk_reset.reset
		.m0_address              (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_003_source0_ready),                                                                           //              cp.ready
		.cp_valid                (burst_adapter_003_source0_valid),                                                                           //                .valid
		.cp_data                 (burst_adapter_003_source0_data),                                                                            //                .data
		.cp_startofpacket        (burst_adapter_003_source0_startofpacket),                                                                   //                .startofpacket
		.cp_endofpacket          (burst_adapter_003_source0_endofpacket),                                                                     //                .endofpacket
		.cp_channel              (burst_adapter_003_source0_channel),                                                                         //                .channel
		.rf_sink_ready           (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (79),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clocks_sys_clk_clk),                                                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                            // clk_reset.reset
		.in_data           (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                                      // (terminated)
		.csr_readdata      (),                                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                      // (terminated)
		.almost_full_data  (),                                                                                                          // (terminated)
		.almost_empty_data (),                                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                                      // (terminated)
		.out_empty         (),                                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                                      // (terminated)
		.out_error         (),                                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                                      // (terminated)
		.out_channel       ()                                                                                                           // (terminated)
	);

	nios_system_addr_router addr_router (
		.sink_ready         (nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_processor_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                 // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                          //       src.ready
		.src_valid          (addr_router_src_valid),                                                                          //          .valid
		.src_data           (addr_router_src_data),                                                                           //          .data
		.src_channel        (addr_router_src_channel),                                                                        //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                                  //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                                     //          .endofpacket
	);

	nios_system_addr_router_001 addr_router_001 (
		.sink_ready         (nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_processor_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                               //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                               //          .valid
		.src_data           (addr_router_001_src_data),                                                                //          .data
		.src_channel        (addr_router_001_src_channel),                                                             //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                       //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                          //          .endofpacket
	);

	nios_system_addr_router_002 addr_router_002 (
		.sink_ready         (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                       // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                                                            //       src.ready
		.src_valid          (addr_router_002_src_valid),                                                                            //          .valid
		.src_data           (addr_router_002_src_data),                                                                             //          .data
		.src_channel        (addr_router_002_src_channel),                                                                          //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                                                    //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                                                       //          .endofpacket
	);

	nios_system_id_router id_router (
		.sink_ready         (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_processor_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                          //       src.ready
		.src_valid          (id_router_src_valid),                                                                          //          .valid
		.src_data           (id_router_src_data),                                                                           //          .data
		.src_channel        (id_router_src_channel),                                                                        //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                                  //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                                     //          .endofpacket
	);

	nios_system_id_router id_router_001 (
		.sink_ready         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                        //       src.ready
		.src_valid          (id_router_001_src_valid),                                                        //          .valid
		.src_data           (id_router_001_src_data),                                                         //          .data
		.src_channel        (id_router_001_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                   //          .endofpacket
	);

	nios_system_id_router_002 id_router_002 (
		.sink_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                             //       src.ready
		.src_valid          (id_router_002_src_valid),                                             //          .valid
		.src_data           (id_router_002_src_data),                                              //          .data
		.src_channel        (id_router_002_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                        //          .endofpacket
	);

	nios_system_id_router_003 id_router_003 (
		.sink_ready         (leds_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (leds_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (leds_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                            //       src.ready
		.src_valid          (id_router_003_src_valid),                                            //          .valid
		.src_data           (id_router_003_src_data),                                             //          .data
		.src_channel        (id_router_003_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                       //          .endofpacket
	);

	nios_system_id_router_003 id_router_004 (
		.sink_ready         (switches_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (switches_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (switches_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (switches_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (switches_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                         // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                //       src.ready
		.src_valid          (id_router_004_src_valid),                                                //          .valid
		.src_data           (id_router_004_src_data),                                                 //          .data
		.src_channel        (id_router_004_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                           //          .endofpacket
	);

	nios_system_id_router_003 id_router_005 (
		.sink_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_005_src_valid),                                                                  //          .valid
		.src_data           (id_router_005_src_data),                                                                   //          .data
		.src_channel        (id_router_005_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                             //          .endofpacket
	);

	nios_system_id_router_006 id_router_006 (
		.sink_ready         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                                     //       src.ready
		.src_valid          (id_router_006_src_valid),                                                                     //          .valid
		.src_data           (id_router_006_src_data),                                                                      //          .data
		.src_channel        (id_router_006_src_channel),                                                                   //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                                             //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                                                //          .endofpacket
	);

	nios_system_id_router_007 id_router_007 (
		.sink_ready         (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                                                   //       src.ready
		.src_valid          (id_router_007_src_valid),                                                                   //          .valid
		.src_data           (id_router_007_src_data),                                                                    //          .data
		.src_channel        (id_router_007_src_channel),                                                                 //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                                           //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                                              //          .endofpacket
	);

	nios_system_id_router_003 id_router_008 (
		.sink_ready         (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                   // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                                                          //       src.ready
		.src_valid          (id_router_008_src_valid),                                                                          //          .valid
		.src_data           (id_router_008_src_data),                                                                           //          .data
		.src_channel        (id_router_008_src_channel),                                                                        //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                                                  //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                                                     //          .endofpacket
	);

	nios_system_id_router_003 id_router_009 (
		.sink_ready         (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (char_drawer_avalon_char_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                   // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                                                          //       src.ready
		.src_valid          (id_router_009_src_valid),                                                                          //          .valid
		.src_data           (id_router_009_src_data),                                                                           //          .data
		.src_channel        (id_router_009_src_channel),                                                                        //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                                                  //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                                                     //          .endofpacket
	);

	nios_system_id_router_006 id_router_010 (
		.sink_ready         (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (char_drawer_avalon_char_buffer_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clocks_sys_clk_clk),                                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                  // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                                                         //       src.ready
		.src_valid          (id_router_010_src_valid),                                                                         //          .valid
		.src_data           (id_router_010_src_data),                                                                          //          .data
		.src_channel        (id_router_010_src_channel),                                                                       //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                                                 //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                                                    //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (94),
		.PKT_DEST_ID_L             (91),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.MAX_OUTSTANDING_RESPONSES (9),
		.PIPELINED                 (0),
		.ST_DATA_W                 (105),
		.ST_CHANNEL_W              (11),
		.VALID_WIDTH               (11),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (clocks_sys_clk_clk),             //       clk.clk
		.reset                  (rst_controller_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_src_data),           //          .data
		.cmd_sink_channel       (addr_router_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (68),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (87),
		.ST_CHANNEL_W              (11),
		.OUT_BYTE_CNT_H            (57),
		.OUT_BURSTWRAP_H           (61),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter (
		.clk                   (clocks_sys_clk_clk),                  //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_002_src_valid),          //     sink0.valid
		.sink0_data            (cmd_xbar_mux_002_src_data),           //          .data
		.sink0_channel         (cmd_xbar_mux_002_src_channel),        //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_002_src_startofpacket),  //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_002_src_endofpacket),    //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_002_src_ready),          //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (59),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURST_SIZE_H          (55),
		.PKT_BURST_SIZE_L          (53),
		.PKT_BURST_TYPE_H          (57),
		.PKT_BURST_TYPE_L          (56),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (78),
		.ST_CHANNEL_W              (11),
		.OUT_BYTE_CNT_H            (47),
		.OUT_BURSTWRAP_H           (52),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_001 (
		.clk                   (clocks_sys_clk_clk),                      //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (width_adapter_002_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_002_src_data),              //          .data
		.sink0_channel         (width_adapter_002_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_002_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_002_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_002_src_ready),             //          .ready
		.source0_valid         (burst_adapter_001_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_001_source0_data),          //          .data
		.source0_channel       (burst_adapter_001_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_001_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_001_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_001_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (68),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (87),
		.ST_CHANNEL_W              (11),
		.OUT_BYTE_CNT_H            (57),
		.OUT_BURSTWRAP_H           (61),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_002 (
		.clk                   (clocks_sys_clk_clk),                      //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_007_src_valid),              //     sink0.valid
		.sink0_data            (cmd_xbar_mux_007_src_data),               //          .data
		.sink0_channel         (cmd_xbar_mux_007_src_channel),            //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_007_src_startofpacket),      //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_007_src_endofpacket),        //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_007_src_ready),              //          .ready
		.source0_valid         (burst_adapter_002_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_002_source0_data),          //          .data
		.source0_channel       (burst_adapter_002_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_002_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_002_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_002_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (59),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURST_SIZE_H          (55),
		.PKT_BURST_SIZE_L          (53),
		.PKT_BURST_TYPE_H          (57),
		.PKT_BURST_TYPE_L          (56),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (78),
		.ST_CHANNEL_W              (11),
		.OUT_BYTE_CNT_H            (47),
		.OUT_BURSTWRAP_H           (52),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_003 (
		.clk                   (clocks_sys_clk_clk),                      //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (width_adapter_004_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_004_src_data),              //          .data
		.sink0_channel         (width_adapter_004_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_004_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_004_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_004_src_ready),             //          .ready
		.source0_valid         (burst_adapter_003_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_003_source0_data),          //          .data
		.source0_channel       (burst_adapter_003_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_003_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_003_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_003_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (nios2_processor_jtag_debug_module_reset_reset), // reset_in0.reset
		.reset_in1  (~reset_reset_n),                                // reset_in1.reset
		.clk        (clocks_sys_clk_clk),                            //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),                // reset_out.reset
		.reset_in2  (1'b0),                                          // (terminated)
		.reset_in3  (1'b0),                                          // (terminated)
		.reset_in4  (1'b0),                                          // (terminated)
		.reset_in5  (1'b0),                                          // (terminated)
		.reset_in6  (1'b0),                                          // (terminated)
		.reset_in7  (1'b0),                                          // (terminated)
		.reset_in8  (1'b0),                                          // (terminated)
		.reset_in9  (1'b0),                                          // (terminated)
		.reset_in10 (1'b0),                                          // (terminated)
		.reset_in11 (1'b0),                                          // (terminated)
		.reset_in12 (1'b0),                                          // (terminated)
		.reset_in13 (1'b0),                                          // (terminated)
		.reset_in14 (1'b0),                                          // (terminated)
		.reset_in15 (1'b0)                                           // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_001 (
		.reset_in0  (~reset_reset_n),                                // reset_in0.reset
		.reset_in1  (nios2_processor_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clk_clk),                                       //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset),            // reset_out.reset
		.reset_in2  (1'b0),                                          // (terminated)
		.reset_in3  (1'b0),                                          // (terminated)
		.reset_in4  (1'b0),                                          // (terminated)
		.reset_in5  (1'b0),                                          // (terminated)
		.reset_in6  (1'b0),                                          // (terminated)
		.reset_in7  (1'b0),                                          // (terminated)
		.reset_in8  (1'b0),                                          // (terminated)
		.reset_in9  (1'b0),                                          // (terminated)
		.reset_in10 (1'b0),                                          // (terminated)
		.reset_in11 (1'b0),                                          // (terminated)
		.reset_in12 (1'b0),                                          // (terminated)
		.reset_in13 (1'b0),                                          // (terminated)
		.reset_in14 (1'b0),                                          // (terminated)
		.reset_in15 (1'b0)                                           // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_002 (
		.reset_in0  (~reset_reset_n),                                // reset_in0.reset
		.reset_in1  (nios2_processor_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clocks_vga_clk_clk),                            //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset),            // reset_out.reset
		.reset_in2  (1'b0),                                          // (terminated)
		.reset_in3  (1'b0),                                          // (terminated)
		.reset_in4  (1'b0),                                          // (terminated)
		.reset_in5  (1'b0),                                          // (terminated)
		.reset_in6  (1'b0),                                          // (terminated)
		.reset_in7  (1'b0),                                          // (terminated)
		.reset_in8  (1'b0),                                          // (terminated)
		.reset_in9  (1'b0),                                          // (terminated)
		.reset_in10 (1'b0),                                          // (terminated)
		.reset_in11 (1'b0),                                          // (terminated)
		.reset_in12 (1'b0),                                          // (terminated)
		.reset_in13 (1'b0),                                          // (terminated)
		.reset_in14 (1'b0),                                          // (terminated)
		.reset_in15 (1'b0)                                           // (terminated)
	);

	nios_system_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clocks_sys_clk_clk),                //        clk.clk
		.reset              (rst_controller_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),           //           .channel
		.sink_data          (limiter_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket)    //           .endofpacket
	);

	nios_system_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                 (clocks_sys_clk_clk),                     //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.sink_ready          (addr_router_001_src_ready),              //      sink.ready
		.sink_channel        (addr_router_001_src_channel),            //          .channel
		.sink_data           (addr_router_001_src_data),               //          .data
		.sink_startofpacket  (addr_router_001_src_startofpacket),      //          .startofpacket
		.sink_endofpacket    (addr_router_001_src_endofpacket),        //          .endofpacket
		.sink_valid          (addr_router_001_src_valid),              //          .valid
		.src0_ready          (cmd_xbar_demux_001_src0_ready),          //      src0.ready
		.src0_valid          (cmd_xbar_demux_001_src0_valid),          //          .valid
		.src0_data           (cmd_xbar_demux_001_src0_data),           //          .data
		.src0_channel        (cmd_xbar_demux_001_src0_channel),        //          .channel
		.src0_startofpacket  (cmd_xbar_demux_001_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_001_src0_endofpacket),    //          .endofpacket
		.src1_ready          (cmd_xbar_demux_001_src1_ready),          //      src1.ready
		.src1_valid          (cmd_xbar_demux_001_src1_valid),          //          .valid
		.src1_data           (cmd_xbar_demux_001_src1_data),           //          .data
		.src1_channel        (cmd_xbar_demux_001_src1_channel),        //          .channel
		.src1_startofpacket  (cmd_xbar_demux_001_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_001_src1_endofpacket),    //          .endofpacket
		.src2_ready          (cmd_xbar_demux_001_src2_ready),          //      src2.ready
		.src2_valid          (cmd_xbar_demux_001_src2_valid),          //          .valid
		.src2_data           (cmd_xbar_demux_001_src2_data),           //          .data
		.src2_channel        (cmd_xbar_demux_001_src2_channel),        //          .channel
		.src2_startofpacket  (cmd_xbar_demux_001_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_001_src2_endofpacket),    //          .endofpacket
		.src3_ready          (cmd_xbar_demux_001_src3_ready),          //      src3.ready
		.src3_valid          (cmd_xbar_demux_001_src3_valid),          //          .valid
		.src3_data           (cmd_xbar_demux_001_src3_data),           //          .data
		.src3_channel        (cmd_xbar_demux_001_src3_channel),        //          .channel
		.src3_startofpacket  (cmd_xbar_demux_001_src3_startofpacket),  //          .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_001_src3_endofpacket),    //          .endofpacket
		.src4_ready          (cmd_xbar_demux_001_src4_ready),          //      src4.ready
		.src4_valid          (cmd_xbar_demux_001_src4_valid),          //          .valid
		.src4_data           (cmd_xbar_demux_001_src4_data),           //          .data
		.src4_channel        (cmd_xbar_demux_001_src4_channel),        //          .channel
		.src4_startofpacket  (cmd_xbar_demux_001_src4_startofpacket),  //          .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_001_src4_endofpacket),    //          .endofpacket
		.src5_ready          (cmd_xbar_demux_001_src5_ready),          //      src5.ready
		.src5_valid          (cmd_xbar_demux_001_src5_valid),          //          .valid
		.src5_data           (cmd_xbar_demux_001_src5_data),           //          .data
		.src5_channel        (cmd_xbar_demux_001_src5_channel),        //          .channel
		.src5_startofpacket  (cmd_xbar_demux_001_src5_startofpacket),  //          .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_001_src5_endofpacket),    //          .endofpacket
		.src6_ready          (cmd_xbar_demux_001_src6_ready),          //      src6.ready
		.src6_valid          (cmd_xbar_demux_001_src6_valid),          //          .valid
		.src6_data           (cmd_xbar_demux_001_src6_data),           //          .data
		.src6_channel        (cmd_xbar_demux_001_src6_channel),        //          .channel
		.src6_startofpacket  (cmd_xbar_demux_001_src6_startofpacket),  //          .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_001_src6_endofpacket),    //          .endofpacket
		.src7_ready          (cmd_xbar_demux_001_src7_ready),          //      src7.ready
		.src7_valid          (cmd_xbar_demux_001_src7_valid),          //          .valid
		.src7_data           (cmd_xbar_demux_001_src7_data),           //          .data
		.src7_channel        (cmd_xbar_demux_001_src7_channel),        //          .channel
		.src7_startofpacket  (cmd_xbar_demux_001_src7_startofpacket),  //          .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_001_src7_endofpacket),    //          .endofpacket
		.src8_ready          (cmd_xbar_demux_001_src8_ready),          //      src8.ready
		.src8_valid          (cmd_xbar_demux_001_src8_valid),          //          .valid
		.src8_data           (cmd_xbar_demux_001_src8_data),           //          .data
		.src8_channel        (cmd_xbar_demux_001_src8_channel),        //          .channel
		.src8_startofpacket  (cmd_xbar_demux_001_src8_startofpacket),  //          .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_001_src8_endofpacket),    //          .endofpacket
		.src9_ready          (cmd_xbar_demux_001_src9_ready),          //      src9.ready
		.src9_valid          (cmd_xbar_demux_001_src9_valid),          //          .valid
		.src9_data           (cmd_xbar_demux_001_src9_data),           //          .data
		.src9_channel        (cmd_xbar_demux_001_src9_channel),        //          .channel
		.src9_startofpacket  (cmd_xbar_demux_001_src9_startofpacket),  //          .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_001_src9_endofpacket),    //          .endofpacket
		.src10_ready         (cmd_xbar_demux_001_src10_ready),         //     src10.ready
		.src10_valid         (cmd_xbar_demux_001_src10_valid),         //          .valid
		.src10_data          (cmd_xbar_demux_001_src10_data),          //          .data
		.src10_channel       (cmd_xbar_demux_001_src10_channel),       //          .channel
		.src10_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //          .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_001_src10_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_002 cmd_xbar_demux_002 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_002_src_ready),             //      sink.ready
		.sink_channel       (addr_router_002_src_channel),           //          .channel
		.sink_data          (addr_router_002_src_data),              //          .data
		.sink_startofpacket (addr_router_002_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_002_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_002_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clocks_sys_clk_clk),                    //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (clocks_sys_clk_clk),                    //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux_002 cmd_xbar_mux_002 (
		.clk                 (clocks_sys_clk_clk),                  //       clk.clk
		.reset               (rst_controller_reset_out_reset),      // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),          //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),          //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),           //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),        //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),  //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),    //          .endofpacket
		.sink0_ready         (width_adapter_src_ready),             //     sink0.ready
		.sink0_valid         (width_adapter_src_valid),             //          .valid
		.sink0_channel       (width_adapter_src_channel),           //          .channel
		.sink0_data          (width_adapter_src_data),              //          .data
		.sink0_startofpacket (width_adapter_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (width_adapter_src_endofpacket),       //          .endofpacket
		.sink1_ready         (width_adapter_001_src_ready),         //     sink1.ready
		.sink1_valid         (width_adapter_001_src_valid),         //          .valid
		.sink1_channel       (width_adapter_001_src_channel),       //          .channel
		.sink1_data          (width_adapter_001_src_data),          //          .data
		.sink1_startofpacket (width_adapter_001_src_startofpacket), //          .startofpacket
		.sink1_endofpacket   (width_adapter_001_src_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux_002 cmd_xbar_mux_007 (
		.clk                 (clocks_sys_clk_clk),                    //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_007_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_007_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_007_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_007_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_007_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_007_src_endofpacket),      //          .endofpacket
		.sink0_ready         (width_adapter_003_src_ready),           //     sink0.ready
		.sink0_valid         (width_adapter_003_src_valid),           //          .valid
		.sink0_channel       (width_adapter_003_src_channel),         //          .channel
		.sink0_data          (width_adapter_003_src_data),            //          .data
		.sink0_startofpacket (width_adapter_003_src_startofpacket),   //          .startofpacket
		.sink0_endofpacket   (width_adapter_003_src_endofpacket),     //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux (
		.clk                (clocks_sys_clk_clk),                //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_002 rsp_xbar_demux_002 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_003 rsp_xbar_demux_003 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_003 rsp_xbar_demux_004 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_003 rsp_xbar_demux_005 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_006 rsp_xbar_demux_006 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_002 rsp_xbar_demux_007 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_007_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_007_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_007_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_007_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_007_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_007_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_003 rsp_xbar_demux_008 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_003 rsp_xbar_demux_009 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_006 rsp_xbar_demux_010 (
		.clk                (clocks_sys_clk_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (clocks_sys_clk_clk),                    //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (width_adapter_005_src_ready),           //     sink2.ready
		.sink2_valid         (width_adapter_005_src_valid),           //          .valid
		.sink2_channel       (width_adapter_005_src_channel),         //          .channel
		.sink2_data          (width_adapter_005_src_data),            //          .data
		.sink2_startofpacket (width_adapter_005_src_startofpacket),   //          .startofpacket
		.sink2_endofpacket   (width_adapter_005_src_endofpacket)      //          .endofpacket
	);

	nios_system_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                  (clocks_sys_clk_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready          (width_adapter_006_src_ready),           //     sink2.ready
		.sink2_valid          (width_adapter_006_src_valid),           //          .valid
		.sink2_channel        (width_adapter_006_src_channel),         //          .channel
		.sink2_data           (width_adapter_006_src_data),            //          .data
		.sink2_startofpacket  (width_adapter_006_src_startofpacket),   //          .startofpacket
		.sink2_endofpacket    (width_adapter_006_src_endofpacket),     //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (width_adapter_007_src_ready),           //     sink6.ready
		.sink6_valid          (width_adapter_007_src_valid),           //          .valid
		.sink6_channel        (width_adapter_007_src_channel),         //          .channel
		.sink6_data           (width_adapter_007_src_data),            //          .data
		.sink6_startofpacket  (width_adapter_007_src_startofpacket),   //          .startofpacket
		.sink6_endofpacket    (width_adapter_007_src_endofpacket),     //          .endofpacket
		.sink7_ready          (width_adapter_008_src_ready),           //     sink7.ready
		.sink7_valid          (width_adapter_008_src_valid),           //          .valid
		.sink7_channel        (width_adapter_008_src_channel),         //          .channel
		.sink7_data           (width_adapter_008_src_data),            //          .data
		.sink7_startofpacket  (width_adapter_008_src_startofpacket),   //          .startofpacket
		.sink7_endofpacket    (width_adapter_008_src_endofpacket),     //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_009_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_009_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (width_adapter_009_src_ready),           //    sink10.ready
		.sink10_valid         (width_adapter_009_src_valid),           //          .valid
		.sink10_channel       (width_adapter_009_src_channel),         //          .channel
		.sink10_data          (width_adapter_009_src_data),            //          .data
		.sink10_startofpacket (width_adapter_009_src_startofpacket),   //          .startofpacket
		.sink10_endofpacket   (width_adapter_009_src_endofpacket)      //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (104),
		.IN_PKT_RESPONSE_STATUS_L      (103),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (105),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (58),
		.OUT_PKT_BYTE_CNT_L            (56),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_PKT_BURST_SIZE_H          (64),
		.OUT_PKT_BURST_SIZE_L          (62),
		.OUT_PKT_RESPONSE_STATUS_H     (86),
		.OUT_PKT_RESPONSE_STATUS_L     (85),
		.OUT_PKT_TRANS_EXCLUSIVE       (55),
		.OUT_PKT_BURST_TYPE_H          (66),
		.OUT_PKT_BURST_TYPE_L          (65),
		.OUT_ST_DATA_W                 (87),
		.ST_CHANNEL_W                  (11),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter (
		.clk                  (clocks_sys_clk_clk),                //       clk.clk
		.reset                (rst_controller_reset_out_reset),    // clk_reset.reset
		.in_valid             (cmd_xbar_demux_src2_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_src2_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_src2_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_src2_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_src2_ready),         //          .ready
		.in_data              (cmd_xbar_demux_src2_data),          //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_src_data),            //          .data
		.out_channel          (width_adapter_src_channel),         //          .channel
		.out_valid            (width_adapter_src_valid),           //          .valid
		.out_ready            (width_adapter_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                             // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (104),
		.IN_PKT_RESPONSE_STATUS_L      (103),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (105),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (58),
		.OUT_PKT_BYTE_CNT_L            (56),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_PKT_BURST_SIZE_H          (64),
		.OUT_PKT_BURST_SIZE_L          (62),
		.OUT_PKT_RESPONSE_STATUS_H     (86),
		.OUT_PKT_RESPONSE_STATUS_L     (85),
		.OUT_PKT_TRANS_EXCLUSIVE       (55),
		.OUT_PKT_BURST_TYPE_H          (66),
		.OUT_PKT_BURST_TYPE_L          (65),
		.OUT_ST_DATA_W                 (87),
		.ST_CHANNEL_W                  (11),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_001 (
		.clk                  (clocks_sys_clk_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src2_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src2_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src2_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src2_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src2_data),          //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_001_src_data),            //          .data
		.out_channel          (width_adapter_001_src_channel),         //          .channel
		.out_valid            (width_adapter_001_src_valid),           //          .valid
		.out_ready            (width_adapter_001_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (104),
		.IN_PKT_RESPONSE_STATUS_L      (103),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (105),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (49),
		.OUT_PKT_BYTE_CNT_L            (47),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_PKT_BURST_SIZE_H          (55),
		.OUT_PKT_BURST_SIZE_L          (53),
		.OUT_PKT_RESPONSE_STATUS_H     (77),
		.OUT_PKT_RESPONSE_STATUS_L     (76),
		.OUT_PKT_TRANS_EXCLUSIVE       (46),
		.OUT_PKT_BURST_TYPE_H          (57),
		.OUT_PKT_BURST_TYPE_L          (56),
		.OUT_ST_DATA_W                 (78),
		.ST_CHANNEL_W                  (11),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_002 (
		.clk                  (clocks_sys_clk_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src6_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src6_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src6_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src6_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src6_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src6_data),          //          .data
		.out_endofpacket      (width_adapter_002_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_002_src_data),            //          .data
		.out_channel          (width_adapter_002_src_channel),         //          .channel
		.out_valid            (width_adapter_002_src_valid),           //          .valid
		.out_ready            (width_adapter_002_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_002_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (104),
		.IN_PKT_RESPONSE_STATUS_L      (103),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (105),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (58),
		.OUT_PKT_BYTE_CNT_L            (56),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_PKT_BURST_SIZE_H          (64),
		.OUT_PKT_BURST_SIZE_L          (62),
		.OUT_PKT_RESPONSE_STATUS_H     (86),
		.OUT_PKT_RESPONSE_STATUS_L     (85),
		.OUT_PKT_TRANS_EXCLUSIVE       (55),
		.OUT_PKT_BURST_TYPE_H          (66),
		.OUT_PKT_BURST_TYPE_L          (65),
		.OUT_ST_DATA_W                 (87),
		.ST_CHANNEL_W                  (11),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_003 (
		.clk                  (clocks_sys_clk_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src7_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src7_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src7_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src7_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src7_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src7_data),          //          .data
		.out_endofpacket      (width_adapter_003_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_003_src_data),            //          .data
		.out_channel          (width_adapter_003_src_channel),         //          .channel
		.out_valid            (width_adapter_003_src_valid),           //          .valid
		.out_ready            (width_adapter_003_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_003_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (104),
		.IN_PKT_RESPONSE_STATUS_L      (103),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (105),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (49),
		.OUT_PKT_BYTE_CNT_L            (47),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_PKT_BURST_SIZE_H          (55),
		.OUT_PKT_BURST_SIZE_L          (53),
		.OUT_PKT_RESPONSE_STATUS_H     (77),
		.OUT_PKT_RESPONSE_STATUS_L     (76),
		.OUT_PKT_TRANS_EXCLUSIVE       (46),
		.OUT_PKT_BURST_TYPE_H          (57),
		.OUT_PKT_BURST_TYPE_L          (56),
		.OUT_ST_DATA_W                 (78),
		.ST_CHANNEL_W                  (11),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_004 (
		.clk                  (clocks_sys_clk_clk),                     //       clk.clk
		.reset                (rst_controller_reset_out_reset),         // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src10_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src10_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src10_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src10_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src10_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src10_data),          //          .data
		.out_endofpacket      (width_adapter_004_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_004_src_data),             //          .data
		.out_channel          (width_adapter_004_src_channel),          //          .channel
		.out_valid            (width_adapter_004_src_valid),            //          .valid
		.out_ready            (width_adapter_004_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_004_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                                  // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (58),
		.IN_PKT_BYTE_CNT_L             (56),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (61),
		.IN_PKT_BURSTWRAP_L            (59),
		.IN_PKT_BURST_SIZE_H           (64),
		.IN_PKT_BURST_SIZE_L           (62),
		.IN_PKT_RESPONSE_STATUS_H      (86),
		.IN_PKT_RESPONSE_STATUS_L      (85),
		.IN_PKT_TRANS_EXCLUSIVE        (55),
		.IN_PKT_BURST_TYPE_H           (66),
		.IN_PKT_BURST_TYPE_L           (65),
		.IN_ST_DATA_W                  (87),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (104),
		.OUT_PKT_RESPONSE_STATUS_L     (103),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (105),
		.ST_CHANNEL_W                  (11),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_005 (
		.clk                  (clocks_sys_clk_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_002_src0_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_002_src0_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_002_src0_ready),         //          .ready
		.in_data              (rsp_xbar_demux_002_src0_data),          //          .data
		.out_endofpacket      (width_adapter_005_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_005_src_data),            //          .data
		.out_channel          (width_adapter_005_src_channel),         //          .channel
		.out_valid            (width_adapter_005_src_valid),           //          .valid
		.out_ready            (width_adapter_005_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_005_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (58),
		.IN_PKT_BYTE_CNT_L             (56),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (61),
		.IN_PKT_BURSTWRAP_L            (59),
		.IN_PKT_BURST_SIZE_H           (64),
		.IN_PKT_BURST_SIZE_L           (62),
		.IN_PKT_RESPONSE_STATUS_H      (86),
		.IN_PKT_RESPONSE_STATUS_L      (85),
		.IN_PKT_TRANS_EXCLUSIVE        (55),
		.IN_PKT_BURST_TYPE_H           (66),
		.IN_PKT_BURST_TYPE_L           (65),
		.IN_ST_DATA_W                  (87),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (104),
		.OUT_PKT_RESPONSE_STATUS_L     (103),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (105),
		.ST_CHANNEL_W                  (11),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_006 (
		.clk                  (clocks_sys_clk_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_002_src1_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_002_src1_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_002_src1_ready),         //          .ready
		.in_data              (rsp_xbar_demux_002_src1_data),          //          .data
		.out_endofpacket      (width_adapter_006_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_006_src_data),            //          .data
		.out_channel          (width_adapter_006_src_channel),         //          .channel
		.out_valid            (width_adapter_006_src_valid),           //          .valid
		.out_ready            (width_adapter_006_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_006_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (49),
		.IN_PKT_BYTE_CNT_L             (47),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (52),
		.IN_PKT_BURSTWRAP_L            (50),
		.IN_PKT_BURST_SIZE_H           (55),
		.IN_PKT_BURST_SIZE_L           (53),
		.IN_PKT_RESPONSE_STATUS_H      (77),
		.IN_PKT_RESPONSE_STATUS_L      (76),
		.IN_PKT_TRANS_EXCLUSIVE        (46),
		.IN_PKT_BURST_TYPE_H           (57),
		.IN_PKT_BURST_TYPE_L           (56),
		.IN_ST_DATA_W                  (78),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (104),
		.OUT_PKT_RESPONSE_STATUS_L     (103),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (105),
		.ST_CHANNEL_W                  (11),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_007 (
		.clk                  (clocks_sys_clk_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_006_src0_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_006_src0_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_006_src0_ready),         //          .ready
		.in_data              (rsp_xbar_demux_006_src0_data),          //          .data
		.out_endofpacket      (width_adapter_007_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_007_src_data),            //          .data
		.out_channel          (width_adapter_007_src_channel),         //          .channel
		.out_valid            (width_adapter_007_src_valid),           //          .valid
		.out_ready            (width_adapter_007_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_007_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (58),
		.IN_PKT_BYTE_CNT_L             (56),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (61),
		.IN_PKT_BURSTWRAP_L            (59),
		.IN_PKT_BURST_SIZE_H           (64),
		.IN_PKT_BURST_SIZE_L           (62),
		.IN_PKT_RESPONSE_STATUS_H      (86),
		.IN_PKT_RESPONSE_STATUS_L      (85),
		.IN_PKT_TRANS_EXCLUSIVE        (55),
		.IN_PKT_BURST_TYPE_H           (66),
		.IN_PKT_BURST_TYPE_L           (65),
		.IN_ST_DATA_W                  (87),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (104),
		.OUT_PKT_RESPONSE_STATUS_L     (103),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (105),
		.ST_CHANNEL_W                  (11),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_008 (
		.clk                  (clocks_sys_clk_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_007_src0_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_007_src0_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_007_src0_ready),         //          .ready
		.in_data              (rsp_xbar_demux_007_src0_data),          //          .data
		.out_endofpacket      (width_adapter_008_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_008_src_data),            //          .data
		.out_channel          (width_adapter_008_src_channel),         //          .channel
		.out_valid            (width_adapter_008_src_valid),           //          .valid
		.out_ready            (width_adapter_008_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_008_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (49),
		.IN_PKT_BYTE_CNT_L             (47),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (52),
		.IN_PKT_BURSTWRAP_L            (50),
		.IN_PKT_BURST_SIZE_H           (55),
		.IN_PKT_BURST_SIZE_L           (53),
		.IN_PKT_RESPONSE_STATUS_H      (77),
		.IN_PKT_RESPONSE_STATUS_L      (76),
		.IN_PKT_TRANS_EXCLUSIVE        (46),
		.IN_PKT_BURST_TYPE_H           (57),
		.IN_PKT_BURST_TYPE_L           (56),
		.IN_ST_DATA_W                  (78),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (104),
		.OUT_PKT_RESPONSE_STATUS_L     (103),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (105),
		.ST_CHANNEL_W                  (11),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_009 (
		.clk                  (clocks_sys_clk_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_010_src0_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_010_src0_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_010_src0_ready),         //          .ready
		.in_data              (rsp_xbar_demux_010_src0_data),          //          .data
		.out_endofpacket      (width_adapter_009_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_009_src_data),            //          .data
		.out_channel          (width_adapter_009_src_channel),         //          .channel
		.out_valid            (width_adapter_009_src_valid),           //          .valid
		.out_ready            (width_adapter_009_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_009_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	nios_system_irq_mapper irq_mapper (
		.clk           (clocks_sys_clk_clk),             //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_processor_d_irq_irq)       //    sender.irq
	);

endmodule
